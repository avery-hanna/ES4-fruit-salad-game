library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ROM is
  port(
	  row : in std_logic_vector(4 downto 0);
	  col : in std_logic_vector(4 downto 0);
	  fruit_color : in std_logic_vector(5 downto 0);
	  clk : in std_logic;
	  color : out std_logic_vector(5 downto 0)
  );
end ROM;

architecture synth of ROM is 
signal address : std_logic_vector(9 downto 0);
begin
	process(clk) is
	begin
		if rising_edge(clk) then
			case address is 

 	 	 	when 0000001101=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000001110=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000001111=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000010000=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000010001=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000101010=> 
 	 	 	 	 <= GFG6FE
 	 	 	when 0000101011=> 
 	 	 	 	 <= GCEBC2
 	 	 	when 0000101100=> 
 	 	 	 	 <= GBD482
 	 	 	when 0000101101=> 
 	 	 	 	 <= G8C460
 	 	 	when 0000101110=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0000101111=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0000110000=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0000110001=> 
 	 	 	 	 <= G8C057
 	 	 	when 0000110010=> 
 	 	 	 	 <= G9CF75
 	 	 	when 0000110011=> 
 	 	 	 	 <= GCE2B0
 	 	 	when 0000110100=> 
 	 	 	 	 <= GEFEE9
 	 	 	when 0000110101=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0001001000=> 
 	 	 	 	 <= GEG0F1
 	 	 	when 0001001001=> 
 	 	 	 	 <= GBD584
 	 	 	when 0001001010=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0001001011=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0001001100=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0001001101=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0001001110=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0001001111=> 
 	 	 	 	 <= G8BG53
 	 	 	when 0001010000=> 
 	 	 	 	 <= G8BF52
 	 	 	when 0001010001=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0001010010=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0001010011=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0001010100=> 
 	 	 	 	 <= G7BD50
 	 	 	when 0001010101=> 
 	 	 	 	 <= G8C869
 	 	 	when 0001010110=> 
 	 	 	 	 <= GDF1D0
 	 	 	when 0001010111=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0001100110=> 
 	 	 	 	 <= GFGEGC
 	 	 	when 0001100111=> 
 	 	 	 	 <= GBE09D
 	 	 	when 0001101000=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0001101001=> 
 	 	 	 	 <= G7BE50
 	 	 	when 0001101010=> 
 	 	 	 	 <= G8BE52
 	 	 	when 0001101011=> 
 	 	 	 	 <= GBD278
 	 	 	when 0001101100=> 
 	 	 	 	 <= GDE99B
 	 	 	when 0001101101=> 
 	 	 	 	 <= GFF9C4
 	 	 	when 0001101110=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0001101111=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0001110000=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0001110001=> 
 	 	 	 	 <= GFFGCF
 	 	 	when 0001110010=> 
 	 	 	 	 <= GEF3BB
 	 	 	when 0001110011=> 
 	 	 	 	 <= GCE08C
 	 	 	when 0001110100=> 
 	 	 	 	 <= G9C862
 	 	 	when 0001110101=> 
 	 	 	 	 <= G8BD50
 	 	 	when 0001110110=> 
 	 	 	 	 <= G7BD50
 	 	 	when 0001110111=> 
 	 	 	 	 <= G9CE73
 	 	 	when 0001111000=> 
 	 	 	 	 <= GFG3F7
 	 	 	when 0010000101=> 
 	 	 	 	 <= GFG8G1
 	 	 	when 0010000110=> 
 	 	 	 	 <= G9CD71
 	 	 	when 0010000111=> 
 	 	 	 	 <= G7BD4G
 	 	 	when 0010001000=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0010001001=> 
 	 	 	 	 <= GCD981
 	 	 	when 0010001010=> 
 	 	 	 	 <= GFFCC9
 	 	 	when 0010001011=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0010001100=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0010001101=> 
 	 	 	 	 <= GFF4CC
 	 	 	when 0010001110=> 
 	 	 	 	 <= GFE6C5
 	 	 	when 0010001111=> 
 	 	 	 	 <= GFE7C6
 	 	 	when 0010010000=> 
 	 	 	 	 <= GFF1CB
 	 	 	when 0010010001=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 0010010010=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0010010011=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0010010100=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0010010101=> 
 	 	 	 	 <= GEF0B5
 	 	 	when 0010010110=> 
 	 	 	 	 <= G9C964
 	 	 	when 0010010111=> 
 	 	 	 	 <= G8BE4G
 	 	 	when 0010011000=> 
 	 	 	 	 <= G8C056
 	 	 	when 0010011001=> 
 	 	 	 	 <= GDF7DE
 	 	 	when 0010011010=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0010100100=> 
 	 	 	 	 <= GFG8G0
 	 	 	when 0010100101=> 
 	 	 	 	 <= G8C767
 	 	 	when 0010100110=> 
 	 	 	 	 <= G8BD50
 	 	 	when 0010100111=> 
 	 	 	 	 <= G8C45D
 	 	 	when 0010101000=> 
 	 	 	 	 <= GEF2BF
 	 	 	when 0010101001=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0010101010=> 
 	 	 	 	 <= GFF9CE
 	 	 	when 0010101011=> 
 	 	 	 	 <= GFD3BF
 	 	 	when 0010101100=> 
 	 	 	 	 <= GFB4B1
 	 	 	when 0010101101=> 
 	 	 	 	 <= GF9G9G
 	 	 	when 0010101110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0010101111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0010110000=> 
 	 	 	 	 <= GF9F9F
 	 	 	when 0010110001=> 
 	 	 	 	 <= GFFBCF
 	 	 	when 0010110010=> 
 	 	 	 	 <= GFB4B1
 	 	 	when 0010110011=> 
 	 	 	 	 <= GFBGB6
 	 	 	when 0010110100=> 
 	 	 	 	 <= GFE3C4
 	 	 	when 0010110101=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0010110110=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0010110111=> 
 	 	 	 	 <= GCDG88
 	 	 	when 0010111000=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0010111001=> 
 	 	 	 	 <= G8BE51
 	 	 	when 0010111010=> 
 	 	 	 	 <= GDF6DC
 	 	 	when 0011000011=> 
 	 	 	 	 <= GFGEGC
 	 	 	when 0011000100=> 
 	 	 	 	 <= G9CD71
 	 	 	when 0011000101=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0011000110=> 
 	 	 	 	 <= G9C862
 	 	 	when 0011000111=> 
 	 	 	 	 <= GFFCC8
 	 	 	when 0011001000=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0011001001=> 
 	 	 	 	 <= GFEBC7
 	 	 	when 0011001010=> 
 	 	 	 	 <= GFB19G
 	 	 	when 0011001011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011001100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011001101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011001110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011001111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011010000=> 
 	 	 	 	 <= GFB4B1
 	 	 	when 0011010001=> 
 	 	 	 	 <= GFEEC9
 	 	 	when 0011010010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011010011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011010100=> 
 	 	 	 	 <= GF9F9F
 	 	 	when 0011010101=> 
 	 	 	 	 <= GFBCB4
 	 	 	when 0011010110=> 
 	 	 	 	 <= GFF1CB
 	 	 	when 0011010111=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0011011000=> 
 	 	 	 	 <= GDEB9C
 	 	 	when 0011011001=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0011011010=> 
 	 	 	 	 <= G8BF54
 	 	 	when 0011011011=> 
 	 	 	 	 <= GEFGEF
 	 	 	when 0011100011=> 
 	 	 	 	 <= GCE19E
 	 	 	when 0011100100=> 
 	 	 	 	 <= G7BD4G
 	 	 	when 0011100101=> 
 	 	 	 	 <= G8C45D
 	 	 	when 0011100110=> 
 	 	 	 	 <= GFFDC8
 	 	 	when 0011100111=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0011101000=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0011101001=> 
 	 	 	 	 <= GFDFC2
 	 	 	when 0011101010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011101011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011101100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011101101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011101110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011101111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011110000=> 
 	 	 	 	 <= GFC0B6
 	 	 	when 0011110001=> 
 	 	 	 	 <= GFE1C3
 	 	 	when 0011110010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011110011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011110100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011110101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0011110110=> 
 	 	 	 	 <= GFB09G
 	 	 	when 0011110111=> 
 	 	 	 	 <= GFECC8
 	 	 	when 0011111000=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 0011111001=> 
 	 	 	 	 <= GDE695
 	 	 	when 0011111010=> 
 	 	 	 	 <= G7BD50
 	 	 	when 0011111011=> 
 	 	 	 	 <= G8C765
 	 	 	when 0011111100=> 
 	 	 	 	 <= GFGDG9
 	 	 	when 0100000010=> 
 	 	 	 	 <= GEG1F2
 	 	 	when 0100000011=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0100000100=> 
 	 	 	 	 <= G7BE50
 	 	 	when 0100000101=> 
 	 	 	 	 <= GEF3BB
 	 	 	when 0100000110=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0100000111=> 
 	 	 	 	 <= GFD0BD
 	 	 	when 0100001000=> 
 	 	 	 	 <= GFB9B3
 	 	 	when 0100001001=> 
 	 	 	 	 <= GFEEC8
 	 	 	when 0100001010=> 
 	 	 	 	 <= GFC8B9
 	 	 	when 0100001011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100001100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100001101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100001110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100001111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100010000=> 
 	 	 	 	 <= GFCEBC
 	 	 	when 0100010001=> 
 	 	 	 	 <= GFD4BF
 	 	 	when 0100010010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100010011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100010100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100010101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100010110=> 
 	 	 	 	 <= GF9G9G
 	 	 	when 0100010111=> 
 	 	 	 	 <= GFD1BE
 	 	 	when 0100011000=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0100011001=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0100011010=> 
 	 	 	 	 <= GBD67B
 	 	 	when 0100011011=> 
 	 	 	 	 <= G7BD50
 	 	 	when 0100011100=> 
 	 	 	 	 <= GCE4B5
 	 	 	when 0100100010=> 
 	 	 	 	 <= GBD687
 	 	 	when 0100100011=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0100100100=> 
 	 	 	 	 <= GBD97G
 	 	 	when 0100100101=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 0100100110=> 
 	 	 	 	 <= GFDBC1
 	 	 	when 0100100111=> 
 	 	 	 	 <= GF9F9G
 	 	 	when 0100101000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100101001=> 
 	 	 	 	 <= GFB3B1
 	 	 	when 0100101010=> 
 	 	 	 	 <= GFF4CC
 	 	 	when 0100101011=> 
 	 	 	 	 <= GFBEB4
 	 	 	when 0100101100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100101101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100101110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100101111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100110000=> 
 	 	 	 	 <= GFDBC1
 	 	 	when 0100110001=> 
 	 	 	 	 <= GFC7B9
 	 	 	when 0100110010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100110011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100110100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0100110101=> 
 	 	 	 	 <= GF9G9G
 	 	 	when 0100110110=> 
 	 	 	 	 <= GFCEBC
 	 	 	when 0100110111=> 
 	 	 	 	 <= GFF5CD
 	 	 	when 0100111000=> 
 	 	 	 	 <= GFDDC1
 	 	 	when 0100111001=> 
 	 	 	 	 <= GFFCCF
 	 	 	when 0100111010=> 
 	 	 	 	 <= GFFECB
 	 	 	when 0100111011=> 
 	 	 	 	 <= G8C056
 	 	 	when 0100111100=> 
 	 	 	 	 <= G8BG56
 	 	 	when 0100111101=> 
 	 	 	 	 <= GFGBG5
 	 	 	when 0101000001=> 
 	 	 	 	 <= GFG7G0
 	 	 	when 0101000010=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0101000011=> 
 	 	 	 	 <= G8BE51
 	 	 	when 0101000100=> 
 	 	 	 	 <= GFFCC8
 	 	 	when 0101000101=> 
 	 	 	 	 <= GFF9CF
 	 	 	when 0101000110=> 
 	 	 	 	 <= GFB09G
 	 	 	when 0101000111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101001000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101001001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101001010=> 
 	 	 	 	 <= GFBBB3
 	 	 	when 0101001011=> 
 	 	 	 	 <= GFF4CD
 	 	 	when 0101001100=> 
 	 	 	 	 <= GFB5B1
 	 	 	when 0101001101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101001110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101001111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101010000=> 
 	 	 	 	 <= GFE7C6
 	 	 	when 0101010001=> 
 	 	 	 	 <= GFBBB3
 	 	 	when 0101010010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101010011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101010100=> 
 	 	 	 	 <= GF9G9G
 	 	 	when 0101010101=> 
 	 	 	 	 <= GFDFC2
 	 	 	when 0101010110=> 
 	 	 	 	 <= GFE7C6
 	 	 	when 0101010111=> 
 	 	 	 	 <= GFB2B0
 	 	 	when 0101011000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101011001=> 
 	 	 	 	 <= GFCBBB
 	 	 	when 0101011010=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0101011011=> 
 	 	 	 	 <= GCDG89
 	 	 	when 0101011100=> 
 	 	 	 	 <= G7BD4G
 	 	 	when 0101011101=> 
 	 	 	 	 <= GCECC3
 	 	 	when 0101100001=> 
 	 	 	 	 <= GCEDC5
 	 	 	when 0101100010=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0101100011=> 
 	 	 	 	 <= GBD273
 	 	 	when 0101100100=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 0101100101=> 
 	 	 	 	 <= GFD5BF
 	 	 	when 0101100110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101100111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101101000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101101001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101101010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101101011=> 
 	 	 	 	 <= GFC5B8
 	 	 	when 0101101100=> 
 	 	 	 	 <= GFEGC9
 	 	 	when 0101101101=> 
 	 	 	 	 <= GFB09G
 	 	 	when 0101101110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101101111=> 
 	 	 	 	 <= GF9G9G
 	 	 	when 0101110000=> 
 	 	 	 	 <= GFF3CC
 	 	 	when 0101110001=> 
 	 	 	 	 <= GFB09G
 	 	 	when 0101110010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101110011=> 
 	 	 	 	 <= GFB5B1
 	 	 	when 0101110100=> 
 	 	 	 	 <= GFEFC9
 	 	 	when 0101110101=> 
 	 	 	 	 <= GFD6BG
 	 	 	when 0101110110=> 
 	 	 	 	 <= GF9G9G
 	 	 	when 0101110111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101111000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0101111001=> 
 	 	 	 	 <= GF9G9G
 	 	 	when 0101111010=> 
 	 	 	 	 <= GFF7CE
 	 	 	when 0101111011=> 
 	 	 	 	 <= GFFCC7
 	 	 	when 0101111100=> 
 	 	 	 	 <= G7BE50
 	 	 	when 0101111101=> 
 	 	 	 	 <= G9CF75
 	 	 	when 0101111110=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0110000001=> 
 	 	 	 	 <= GBD686
 	 	 	when 0110000010=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0110000011=> 
 	 	 	 	 <= GDE898
 	 	 	when 0110000100=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0110000101=> 
 	 	 	 	 <= GFCFBD
 	 	 	when 0110000110=> 
 	 	 	 	 <= GF9G9G
 	 	 	when 0110000111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0110001000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0110001001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0110001010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0110001011=> 
 	 	 	 	 <= GG9G9F
 	 	 	when 0110001100=> 
 	 	 	 	 <= GFD3BF
 	 	 	when 0110001101=> 
 	 	 	 	 <= GFE3C5
 	 	 	when 0110001110=> 
 	 	 	 	 <= GF9F9G
 	 	 	when 0110001111=> 
 	 	 	 	 <= GF9G9G
 	 	 	when 0110010000=> 
 	 	 	 	 <= GFF6CD
 	 	 	when 0110010001=> 
 	 	 	 	 <= GF9F9F
 	 	 	when 0110010010=> 
 	 	 	 	 <= GFBGB5
 	 	 	when 0110010011=> 
 	 	 	 	 <= GFF5CD
 	 	 	when 0110010100=> 
 	 	 	 	 <= GFC5B8
 	 	 	when 0110010101=> 
 	 	 	 	 <= GF9F9F
 	 	 	when 0110010110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0110010111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0110011000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0110011001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0110011010=> 
 	 	 	 	 <= GFD9C0
 	 	 	when 0110011011=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 0110011100=> 
 	 	 	 	 <= G9CB66
 	 	 	when 0110011101=> 
 	 	 	 	 <= G8BE51
 	 	 	when 0110011110=> 
 	 	 	 	 <= GFGDGB
 	 	 	when 0110100000=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0110100001=> 
 	 	 	 	 <= G8C664
 	 	 	when 0110100010=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0110100011=> 
 	 	 	 	 <= GFF8C3
 	 	 	when 0110100100=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0110100101=> 
 	 	 	 	 <= GFF9CF
 	 	 	when 0110100110=> 
 	 	 	 	 <= GFD9C0
 	 	 	when 0110100111=> 
 	 	 	 	 <= GFC7B9
 	 	 	when 0110101000=> 
 	 	 	 	 <= GFBCB4
 	 	 	when 0110101001=> 
 	 	 	 	 <= GFB09G
 	 	 	when 0110101010=> 
 	 	 	 	 <= GF9F9G
 	 	 	when 0110101011=> 
 	 	 	 	 <= GF9F9F
 	 	 	when 0110101100=> 
 	 	 	 	 <= GF9F9F
 	 	 	when 0110101101=> 
 	 	 	 	 <= GFE1C4
 	 	 	when 0110101110=> 
 	 	 	 	 <= GFD9C0
 	 	 	when 0110101111=> 
 	 	 	 	 <= GFC1B6
 	 	 	when 0110110000=> 
 	 	 	 	 <= GFEDC8
 	 	 	when 0110110001=> 
 	 	 	 	 <= GFCFBD
 	 	 	when 0110110010=> 
 	 	 	 	 <= GFF2CC
 	 	 	when 0110110011=> 
 	 	 	 	 <= GFB9B3
 	 	 	when 0110110100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0110110101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0110110110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0110110111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0110111000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0110111001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0110111010=> 
 	 	 	 	 <= GFC2B7
 	 	 	when 0110111011=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 0110111100=> 
 	 	 	 	 <= GBDB80
 	 	 	when 0110111101=> 
 	 	 	 	 <= G8BD4G
 	 	 	when 0110111110=> 
 	 	 	 	 <= GEFGEE
 	 	 	when 0111000000=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0111000001=> 
 	 	 	 	 <= G8BE51
 	 	 	when 0111000010=> 
 	 	 	 	 <= G7BD50
 	 	 	when 0111000011=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0111000100=> 
 	 	 	 	 <= GFFGD0
 	 	 	when 0111000101=> 
 	 	 	 	 <= GFD5BF
 	 	 	when 0111000110=> 
 	 	 	 	 <= GFD2BE
 	 	 	when 0111000111=> 
 	 	 	 	 <= GFDBC0
 	 	 	when 0111001000=> 
 	 	 	 	 <= GFE7C6
 	 	 	when 0111001001=> 
 	 	 	 	 <= GFF3CC
 	 	 	when 0111001010=> 
 	 	 	 	 <= GFF6CD
 	 	 	when 0111001011=> 
 	 	 	 	 <= GFECC8
 	 	 	when 0111001100=> 
 	 	 	 	 <= GFDFC2
 	 	 	when 0111001101=> 
 	 	 	 	 <= GFE1C3
 	 	 	when 0111001110=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0111001111=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 0111010000=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0111010001=> 
 	 	 	 	 <= GFE8C6
 	 	 	when 0111010010=> 
 	 	 	 	 <= GFB1B0
 	 	 	when 0111010011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0111010100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0111010101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0111010110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0111010111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0111011000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0111011001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0111011010=> 
 	 	 	 	 <= GFB4B1
 	 	 	when 0111011011=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0111011100=> 
 	 	 	 	 <= GDE491
 	 	 	when 0111011101=> 
 	 	 	 	 <= G8BD50
 	 	 	when 0111011110=> 
 	 	 	 	 <= GDF5D9
 	 	 	when 0111100000=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0111100001=> 
 	 	 	 	 <= G8BD50
 	 	 	when 0111100010=> 
 	 	 	 	 <= G8BE51
 	 	 	when 0111100011=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0111100100=> 
 	 	 	 	 <= GFE6C6
 	 	 	when 0111100101=> 
 	 	 	 	 <= GF9F9F
 	 	 	when 0111100110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0111100111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0111101000=> 
 	 	 	 	 <= GF9G9F
 	 	 	when 0111101001=> 
 	 	 	 	 <= GF9F9F
 	 	 	when 0111101010=> 
 	 	 	 	 <= GF9F9G
 	 	 	when 0111101011=> 
 	 	 	 	 <= GFB6B2
 	 	 	when 0111101100=> 
 	 	 	 	 <= GFC3B7
 	 	 	when 0111101101=> 
 	 	 	 	 <= GFE2C4
 	 	 	when 0111101110=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0111101111=> 
 	 	 	 	 <= GGG0D0
 	 	 	when 0111110000=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0111110001=> 
 	 	 	 	 <= GFF8CE
 	 	 	when 0111110010=> 
 	 	 	 	 <= GFE8C7
 	 	 	when 0111110011=> 
 	 	 	 	 <= GFDDC1
 	 	 	when 0111110100=> 
 	 	 	 	 <= GFCGBD
 	 	 	when 0111110101=> 
 	 	 	 	 <= GFC2B7
 	 	 	when 0111110110=> 
 	 	 	 	 <= GFB5B1
 	 	 	when 0111110111=> 
 	 	 	 	 <= GF9F9F
 	 	 	when 0111111000=> 
 	 	 	 	 <= GG9F9G
 	 	 	when 0111111001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 0111111010=> 
 	 	 	 	 <= GFBDB4
 	 	 	when 0111111011=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0111111100=> 
 	 	 	 	 <= GDE797
 	 	 	when 0111111101=> 
 	 	 	 	 <= G8BE50
 	 	 	when 0111111110=> 
 	 	 	 	 <= GDF2D2
 	 	 	when 1000000000=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1000000001=> 
 	 	 	 	 <= G8BE50
 	 	 	when 1000000010=> 
 	 	 	 	 <= G8BE50
 	 	 	when 1000000011=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1000000100=> 
 	 	 	 	 <= GFE3C4
 	 	 	when 1000000101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1000000110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1000000111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1000001000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1000001001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1000001010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1000001011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1000001100=> 
 	 	 	 	 <= GG9F9G
 	 	 	when 1000001101=> 
 	 	 	 	 <= GFCGBD
 	 	 	when 1000001110=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1000001111=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1000010000=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1000010001=> 
 	 	 	 	 <= GFC0B6
 	 	 	when 1000010010=> 
 	 	 	 	 <= GFB9B3
 	 	 	when 1000010011=> 
 	 	 	 	 <= GFC5B8
 	 	 	when 1000010100=> 
 	 	 	 	 <= GFD2BE
 	 	 	when 1000010101=> 
 	 	 	 	 <= GFDGC3
 	 	 	when 1000010110=> 
 	 	 	 	 <= GFEDC8
 	 	 	when 1000010111=> 
 	 	 	 	 <= GFF7CD
 	 	 	when 1000011000=> 
 	 	 	 	 <= GFF2CC
 	 	 	when 1000011001=> 
 	 	 	 	 <= GFE6C5
 	 	 	when 1000011010=> 
 	 	 	 	 <= GFE9C7
 	 	 	when 1000011011=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1000011100=> 
 	 	 	 	 <= GCE390
 	 	 	when 1000011101=> 
 	 	 	 	 <= G8BE50
 	 	 	when 1000011110=> 
 	 	 	 	 <= GDF4D6
 	 	 	when 1000100000=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1000100001=> 
 	 	 	 	 <= G8C25D
 	 	 	when 1000100010=> 
 	 	 	 	 <= G8BE50
 	 	 	when 1000100011=> 
 	 	 	 	 <= GFFFCE
 	 	 	when 1000100100=> 
 	 	 	 	 <= GFEDC8
 	 	 	when 1000100101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1000100110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1000100111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1000101000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1000101001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1000101010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1000101011=> 
 	 	 	 	 <= GG9G9F
 	 	 	when 1000101100=> 
 	 	 	 	 <= GFCGBD
 	 	 	when 1000101101=> 
 	 	 	 	 <= GFF2CB
 	 	 	when 1000101110=> 
 	 	 	 	 <= GFB8B3
 	 	 	when 1000101111=> 
 	 	 	 	 <= GFF5CD
 	 	 	when 1000110000=> 
 	 	 	 	 <= GFF0CB
 	 	 	when 1000110001=> 
 	 	 	 	 <= GFEFC9
 	 	 	when 1000110010=> 
 	 	 	 	 <= GFB09G
 	 	 	when 1000110011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1000110100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1000110101=> 
 	 	 	 	 <= GF9F9G
 	 	 	when 1000110110=> 
 	 	 	 	 <= GG9F9G
 	 	 	when 1000110111=> 
 	 	 	 	 <= GG9F9G
 	 	 	when 1000111000=> 
 	 	 	 	 <= GFB09G
 	 	 	when 1000111001=> 
 	 	 	 	 <= GFBDB4
 	 	 	when 1000111010=> 
 	 	 	 	 <= GFEBC7
 	 	 	when 1000111011=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1000111100=> 
 	 	 	 	 <= GCDF87
 	 	 	when 1000111101=> 
 	 	 	 	 <= G7BD4G
 	 	 	when 1000111110=> 
 	 	 	 	 <= GEFCE6
 	 	 	when 1001000001=> 
 	 	 	 	 <= G9D17B
 	 	 	when 1001000010=> 
 	 	 	 	 <= G8BE50
 	 	 	when 1001000011=> 
 	 	 	 	 <= GEF2B8
 	 	 	when 1001000100=> 
 	 	 	 	 <= GFFDCG
 	 	 	when 1001000101=> 
 	 	 	 	 <= GF9G9G
 	 	 	when 1001000110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001000111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001001000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001001001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001001010=> 
 	 	 	 	 <= GFB09G
 	 	 	when 1001001011=> 
 	 	 	 	 <= GFE1C3
 	 	 	when 1001001100=> 
 	 	 	 	 <= GFE5C5
 	 	 	when 1001001101=> 
 	 	 	 	 <= GFB1B0
 	 	 	when 1001001110=> 
 	 	 	 	 <= GF9F9F
 	 	 	when 1001001111=> 
 	 	 	 	 <= GFF5CD
 	 	 	when 1001010000=> 
 	 	 	 	 <= GF9G9G
 	 	 	when 1001010001=> 
 	 	 	 	 <= GFD4BF
 	 	 	when 1001010010=> 
 	 	 	 	 <= GFE2C4
 	 	 	when 1001010011=> 
 	 	 	 	 <= GF9F9F
 	 	 	when 1001010100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001010101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001010110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001010111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001011000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001011001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001011010=> 
 	 	 	 	 <= GFD0BD
 	 	 	when 1001011011=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1001011100=> 
 	 	 	 	 <= GBD378
 	 	 	when 1001011101=> 
 	 	 	 	 <= G7BD50
 	 	 	when 1001011110=> 
 	 	 	 	 <= GFG9G3
 	 	 	when 1001100001=> 
 	 	 	 	 <= GCE5B6
 	 	 	when 1001100010=> 
 	 	 	 	 <= G8BE50
 	 	 	when 1001100011=> 
 	 	 	 	 <= GCDG89
 	 	 	when 1001100100=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1001100101=> 
 	 	 	 	 <= GFC1B6
 	 	 	when 1001100110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001100111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001101000=> 
 	 	 	 	 <= GF9F9F
 	 	 	when 1001101001=> 
 	 	 	 	 <= GFB6B2
 	 	 	when 1001101010=> 
 	 	 	 	 <= GFF0C9
 	 	 	when 1001101011=> 
 	 	 	 	 <= GFD3BF
 	 	 	when 1001101100=> 
 	 	 	 	 <= GF9F9G
 	 	 	when 1001101101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001101110=> 
 	 	 	 	 <= GF9G9G
 	 	 	when 1001101111=> 
 	 	 	 	 <= GFF4CD
 	 	 	when 1001110000=> 
 	 	 	 	 <= GF9F9G
 	 	 	when 1001110001=> 
 	 	 	 	 <= GF9F9G
 	 	 	when 1001110010=> 
 	 	 	 	 <= GFE2C4
 	 	 	when 1001110011=> 
 	 	 	 	 <= GFD3BF
 	 	 	when 1001110100=> 
 	 	 	 	 <= GG9F9G
 	 	 	when 1001110101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001110110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001110111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001111000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1001111001=> 
 	 	 	 	 <= GG9F9G
 	 	 	when 1001111010=> 
 	 	 	 	 <= GFE6C5
 	 	 	when 1001111011=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1001111100=> 
 	 	 	 	 <= G8C15B
 	 	 	when 1001111101=> 
 	 	 	 	 <= G8C766
 	 	 	when 1001111110=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1010000001=> 
 	 	 	 	 <= GEG0EG
 	 	 	when 1010000010=> 
 	 	 	 	 <= G7BD50
 	 	 	when 1010000011=> 
 	 	 	 	 <= G8C660
 	 	 	when 1010000100=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1010000101=> 
 	 	 	 	 <= GFE5C5
 	 	 	when 1010000110=> 
 	 	 	 	 <= GF9F9F
 	 	 	when 1010000111=> 
 	 	 	 	 <= GG9F9G
 	 	 	when 1010001000=> 
 	 	 	 	 <= GFC1B6
 	 	 	when 1010001001=> 
 	 	 	 	 <= GFF5CD
 	 	 	when 1010001010=> 
 	 	 	 	 <= GFC3B7
 	 	 	when 1010001011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1010001100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1010001101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1010001110=> 
 	 	 	 	 <= GFB9B3
 	 	 	when 1010001111=> 
 	 	 	 	 <= GFE8C6
 	 	 	when 1010010000=> 
 	 	 	 	 <= GF9F9G
 	 	 	when 1010010001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1010010010=> 
 	 	 	 	 <= GFB09G
 	 	 	when 1010010011=> 
 	 	 	 	 <= GFEFC9
 	 	 	when 1010010100=> 
 	 	 	 	 <= GFC6B8
 	 	 	when 1010010101=> 
 	 	 	 	 <= GG9F9F
 	 	 	when 1010010110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1010010111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1010011000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1010011001=> 
 	 	 	 	 <= GFB5B1
 	 	 	when 1010011010=> 
 	 	 	 	 <= GFFGD0
 	 	 	when 1010011011=> 
 	 	 	 	 <= GEEFB3
 	 	 	when 1010011100=> 
 	 	 	 	 <= G7BD4G
 	 	 	when 1010011101=> 
 	 	 	 	 <= GCE29G
 	 	 	when 1010100001=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1010100010=> 
 	 	 	 	 <= G9CC6G
 	 	 	when 1010100011=> 
 	 	 	 	 <= G8BD50
 	 	 	when 1010100100=> 
 	 	 	 	 <= GDEEB0
 	 	 	when 1010100101=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1010100110=> 
 	 	 	 	 <= GFE0C3
 	 	 	when 1010100111=> 
 	 	 	 	 <= GFD3BF
 	 	 	when 1010101000=> 
 	 	 	 	 <= GFF1CB
 	 	 	when 1010101001=> 
 	 	 	 	 <= GFB7B2
 	 	 	when 1010101010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1010101011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1010101100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1010101101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1010101110=> 
 	 	 	 	 <= GFC6B8
 	 	 	when 1010101111=> 
 	 	 	 	 <= GFDCC1
 	 	 	when 1010110000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1010110001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1010110010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1010110011=> 
 	 	 	 	 <= GFB5B1
 	 	 	when 1010110100=> 
 	 	 	 	 <= GFF4CC
 	 	 	when 1010110101=> 
 	 	 	 	 <= GFBCB4
 	 	 	when 1010110110=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1010110111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1010111000=> 
 	 	 	 	 <= GF9G9F
 	 	 	when 1010111001=> 
 	 	 	 	 <= GFE0C3
 	 	 	when 1010111010=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1010111011=> 
 	 	 	 	 <= G9CG70
 	 	 	when 1010111100=> 
 	 	 	 	 <= G8BE50
 	 	 	when 1010111101=> 
 	 	 	 	 <= GEG3F6
 	 	 	when 1011000010=> 
 	 	 	 	 <= GDF5D8
 	 	 	when 1011000011=> 
 	 	 	 	 <= G7BD50
 	 	 	when 1011000100=> 
 	 	 	 	 <= G8C65G
 	 	 	when 1011000101=> 
 	 	 	 	 <= GFFGCF
 	 	 	when 1011000110=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1011000111=> 
 	 	 	 	 <= GFF0CB
 	 	 	when 1011001000=> 
 	 	 	 	 <= GFB19G
 	 	 	when 1011001001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011001010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011001011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011001100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011001101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011001110=> 
 	 	 	 	 <= GFD3BF
 	 	 	when 1011001111=> 
 	 	 	 	 <= GFCFBD
 	 	 	when 1011010000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011010001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011010010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011010011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011010100=> 
 	 	 	 	 <= GFBDB4
 	 	 	when 1011010101=> 
 	 	 	 	 <= GFF4CC
 	 	 	when 1011010110=> 
 	 	 	 	 <= GFB4B1
 	 	 	when 1011010111=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011011000=> 
 	 	 	 	 <= GFC4B8
 	 	 	when 1011011001=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1011011010=> 
 	 	 	 	 <= GEF0B5
 	 	 	when 1011011011=> 
 	 	 	 	 <= G7BD4G
 	 	 	when 1011011100=> 
 	 	 	 	 <= GBD687
 	 	 	when 1011011101=> 
 	 	 	 	 <= GFGFGG
 	 	 	when 1011100010=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1011100011=> 
 	 	 	 	 <= G9D07B
 	 	 	when 1011100100=> 
 	 	 	 	 <= G7BE50
 	 	 	when 1011100101=> 
 	 	 	 	 <= GBDB80
 	 	 	when 1011100110=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1011100111=> 
 	 	 	 	 <= GFF7CE
 	 	 	when 1011101000=> 
 	 	 	 	 <= GFB09G
 	 	 	when 1011101001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011101010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011101011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011101100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011101101=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011101110=> 
 	 	 	 	 <= GFE0C3
 	 	 	when 1011101111=> 
 	 	 	 	 <= GFC2B6
 	 	 	when 1011110000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011110001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011110010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011110011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1011110100=> 
 	 	 	 	 <= GF9G9G
 	 	 	when 1011110101=> 
 	 	 	 	 <= GFC7B9
 	 	 	when 1011110110=> 
 	 	 	 	 <= GFEFC9
 	 	 	when 1011110111=> 
 	 	 	 	 <= GFD0BD
 	 	 	when 1011111000=> 
 	 	 	 	 <= GFFDCG
 	 	 	when 1011111001=> 
 	 	 	 	 <= GFFECC
 	 	 	when 1011111010=> 
 	 	 	 	 <= G8C45D
 	 	 	when 1011111011=> 
 	 	 	 	 <= G8BG54
 	 	 	when 1011111100=> 
 	 	 	 	 <= GFG5FB
 	 	 	when 1100000011=> 
 	 	 	 	 <= GFG6FD
 	 	 	when 1100000100=> 
 	 	 	 	 <= G8C15B
 	 	 	when 1100000101=> 
 	 	 	 	 <= G7BD50
 	 	 	when 1100000110=> 
 	 	 	 	 <= GDE798
 	 	 	when 1100000111=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1100001000=> 
 	 	 	 	 <= GFEDC8
 	 	 	when 1100001001=> 
 	 	 	 	 <= GFB3B1
 	 	 	when 1100001010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1100001011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1100001100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1100001101=> 
 	 	 	 	 <= GF9G9F
 	 	 	when 1100001110=> 
 	 	 	 	 <= GFEDC8
 	 	 	when 1100001111=> 
 	 	 	 	 <= GFB5B1
 	 	 	when 1100010000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1100010001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1100010010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1100010011=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1100010100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1100010101=> 
 	 	 	 	 <= GF9F9F
 	 	 	when 1100010110=> 
 	 	 	 	 <= GFF0CB
 	 	 	when 1100010111=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1100011000=> 
 	 	 	 	 <= GFFGCF
 	 	 	when 1100011001=> 
 	 	 	 	 <= G9CE6C
 	 	 	when 1100011010=> 
 	 	 	 	 <= G7BD4G
 	 	 	when 1100011011=> 
 	 	 	 	 <= GDEFCB
 	 	 	when 1100011100=> 
 	 	 	 	 <= GGGFGG
 	 	 	when 1100100100=> 
 	 	 	 	 <= GEFCE6
 	 	 	when 1100100101=> 
 	 	 	 	 <= G8BF53
 	 	 	when 1100100110=> 
 	 	 	 	 <= G8BE50
 	 	 	when 1100100111=> 
 	 	 	 	 <= GDE391
 	 	 	when 1100101000=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 1100101001=> 
 	 	 	 	 <= GFFBCF
 	 	 	when 1100101010=> 
 	 	 	 	 <= GFCDBC
 	 	 	when 1100101011=> 
 	 	 	 	 <= GF9G9G
 	 	 	when 1100101100=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1100101101=> 
 	 	 	 	 <= GF9F9F
 	 	 	when 1100101110=> 
 	 	 	 	 <= GFF7CE
 	 	 	when 1100101111=> 
 	 	 	 	 <= GF9F9F
 	 	 	when 1100110000=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1100110001=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1100110010=> 
 	 	 	 	 <= GG9G9G
 	 	 	when 1100110011=> 
 	 	 	 	 <= GF9G9G
 	 	 	when 1100110100=> 
 	 	 	 	 <= GFB6B1
 	 	 	when 1100110101=> 
 	 	 	 	 <= GFE1C3
 	 	 	when 1100110110=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1100110111=> 
 	 	 	 	 <= GFFECB
 	 	 	when 1100111000=> 
 	 	 	 	 <= G9CD6B
 	 	 	when 1100111001=> 
 	 	 	 	 <= G8BD50
 	 	 	when 1100111010=> 
 	 	 	 	 <= GBDG9B
 	 	 	when 1100111011=> 
 	 	 	 	 <= GGGFGF
 	 	 	when 1101000100=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1101000101=> 
 	 	 	 	 <= GEF9E1
 	 	 	when 1101000110=> 
 	 	 	 	 <= G8BG56
 	 	 	when 1101000111=> 
 	 	 	 	 <= G8BD4G
 	 	 	when 1101001000=> 
 	 	 	 	 <= GBD478
 	 	 	when 1101001001=> 
 	 	 	 	 <= GFFDC9
 	 	 	when 1101001010=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1101001011=> 
 	 	 	 	 <= GFF8CE
 	 	 	when 1101001100=> 
 	 	 	 	 <= GFDBC1
 	 	 	when 1101001101=> 
 	 	 	 	 <= GFD2BE
 	 	 	when 1101001110=> 
 	 	 	 	 <= GFFFD0
 	 	 	when 1101001111=> 
 	 	 	 	 <= GFC5B8
 	 	 	when 1101010000=> 
 	 	 	 	 <= GFB5B1
 	 	 	when 1101010001=> 
 	 	 	 	 <= GFBDB4
 	 	 	when 1101010010=> 
 	 	 	 	 <= GFCDBC
 	 	 	when 1101010011=> 
 	 	 	 	 <= GFE6C6
 	 	 	when 1101010100=> 
 	 	 	 	 <= GFFGD0
 	 	 	when 1101010101=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 1101010110=> 
 	 	 	 	 <= GEEGB4
 	 	 	when 1101010111=> 
 	 	 	 	 <= G8C45D
 	 	 	when 1101011000=> 
 	 	 	 	 <= G8BD4G
 	 	 	when 1101011001=> 
 	 	 	 	 <= GBE09E
 	 	 	when 1101011010=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1101100110=> 
 	 	 	 	 <= GEG2F3
 	 	 	when 1101100111=> 
 	 	 	 	 <= G9C96C
 	 	 	when 1101101000=> 
 	 	 	 	 <= G8BD50
 	 	 	when 1101101001=> 
 	 	 	 	 <= G8C055
 	 	 	when 1101101010=> 
 	 	 	 	 <= GCDE87
 	 	 	when 1101101011=> 
 	 	 	 	 <= GFFBC5
 	 	 	when 1101101100=> 
 	 	 	 	 <= GGG0D1
 	 	 	when 1101101101=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 1101101110=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1101101111=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1101110000=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1101110001=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1101110010=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1101110011=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1101110100=> 
 	 	 	 	 <= GEEGB4
 	 	 	when 1101110101=> 
 	 	 	 	 <= G9CG6G
 	 	 	when 1101110110=> 
 	 	 	 	 <= G8BD50
 	 	 	when 1101110111=> 
 	 	 	 	 <= G8BG55
 	 	 	when 1101111000=> 
 	 	 	 	 <= GDEGCC
 	 	 	when 1101111001=> 
 	 	 	 	 <= GGGFGG
 	 	 	when 1110000111=> 
 	 	 	 	 <= GFGEGD
 	 	 	when 1110001000=> 
 	 	 	 	 <= GCE8BD
 	 	 	when 1110001001=> 
 	 	 	 	 <= G8C159
 	 	 	when 1110001010=> 
 	 	 	 	 <= G8BD50
 	 	 	when 1110001011=> 
 	 	 	 	 <= G8BE50
 	 	 	when 1110001100=> 
 	 	 	 	 <= G9C864
 	 	 	when 1110001101=> 
 	 	 	 	 <= GCD881
 	 	 	when 1110001110=> 
 	 	 	 	 <= GCE38G
 	 	 	when 1110001111=> 
 	 	 	 	 <= GDE796
 	 	 	when 1110010000=> 
 	 	 	 	 <= GDE694
 	 	 	when 1110010001=> 
 	 	 	 	 <= GCDG89
 	 	 	when 1110010010=> 
 	 	 	 	 <= GBD374
 	 	 	when 1110010011=> 
 	 	 	 	 <= G8C157
 	 	 	when 1110010100=> 
 	 	 	 	 <= G7BD50
 	 	 	when 1110010101=> 
 	 	 	 	 <= G8BE50
 	 	 	when 1110010110=> 
 	 	 	 	 <= GBD889
 	 	 	when 1110010111=> 
 	 	 	 	 <= GFG5FC
 	 	 	when 1110011000=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1110101001=> 
 	 	 	 	 <= GFGDG8
 	 	 	when 1110101010=> 
 	 	 	 	 <= GDEFCB
 	 	 	when 1110101011=> 
 	 	 	 	 <= G9D17C
 	 	 	when 1110101100=> 
 	 	 	 	 <= G8BF53
 	 	 	when 1110101101=> 
 	 	 	 	 <= G8BD50
 	 	 	when 1110101110=> 
 	 	 	 	 <= G8BE50
 	 	 	when 1110101111=> 
 	 	 	 	 <= G8BE50
 	 	 	when 1110110000=> 
 	 	 	 	 <= G8BE50
 	 	 	when 1110110001=> 
 	 	 	 	 <= G8BD50
 	 	 	when 1110110010=> 
 	 	 	 	 <= G8BE4G
 	 	 	when 1110110011=> 
 	 	 	 	 <= G9C869
 	 	 	when 1110110100=> 
 	 	 	 	 <= GCE3B2
 	 	 	when 1110110101=> 
 	 	 	 	 <= GFG4F8
 	 	 	when 1110110110=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1111001011=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1111001100=> 
 	 	 	 	 <= GFGFGE
 	 	 	when 1111001101=> 
 	 	 	 	 <= GEG2F3
 	 	 	when 1111001110=> 
 	 	 	 	 <= GEF8DF
 	 	 	when 1111001111=> 
 	 	 	 	 <= GDF5D7
 	 	 	when 1111010000=> 
 	 	 	 	 <= GDF6DB
 	 	 	when 1111010001=> 
 	 	 	 	 <= GEFEEB
 	 	 	when 1111010010=> 
 	 	 	 	 <= GFGCG6
 	 	 	when 1111010011=> 
 	 	 	 	 <= GFGFGF 
 	 	 end case; 
     	 end if;  
     end process; 
 address <= row & col; 
 end;