library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ROM is
  port(
	  row : in std_logic_vector(7 downto 0);
	  col : in std_logic_vector(7 downto 0);
	  fruit_color : in std_logic_vector(5 downto 0);
	  clk : in std_logic;
	  color : out std_logic_vector(5 downto 0)
  );
end ROM;

architecture synth of ROM is 
signal address : std_logic_vector(9 downto 0);
begin
	process(clk) is
	begin
		if rising_edge(clk) then
			case address is 

 	 	 	when "0000001101000010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000001101000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000001101000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000001101000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000001101000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000001101000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000010001000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010001000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010001000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010001000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010001000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010001000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010001000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010001000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010001001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010001001001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000010100111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010101000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010101000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010101000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010101000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010101000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010101000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010101000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010101000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010101001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010101001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010101001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011000111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011000111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011001000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011001000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011001000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011001000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011001000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011001000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011001000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011001000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011001001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011001001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011001001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011001001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011100111110" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000011100111111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000011101000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011101000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011101000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011101000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011101000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011101000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011101000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011101000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011101001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011101001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011101001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011101001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011101001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100000111101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000100000111110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000100000111111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000100001000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100001000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100001000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100001000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100001000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100001000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100001000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100001000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100001001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100001001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100001001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100001001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100001001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100100111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100100111111" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000100101000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100101000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100101000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100101000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100101000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100101000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100101000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100101000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100101001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100101001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100101001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100101001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100101001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100101001101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101000111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101000111111" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000101001000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101001000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101001000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101001000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101001000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101001000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101001000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101001000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101001001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101001001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101001001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101001001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101001001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101001001101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101100111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101100111111" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000101101000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101101000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101101000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101101000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101101000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101101000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101101000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101101000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101101001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101101001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101101001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101101001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101101001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101101001101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110000111101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000110000111110" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0000110000111111" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000110001000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110001000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110001000010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0000110001000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110001000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110001000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110001000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110001000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110001001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110001001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110001001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110001001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110001001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110001001101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110100101000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000110100101010" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000110100101011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000110100101100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000110100101101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0000110100111001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0000110100111010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000110100111011" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000110100111100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000110100111110" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0000110100111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110101000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110101000001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000110101000010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000110101000011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000110101000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110101000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110101000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110101000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110101001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110101001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110101001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110101001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110101001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110101001101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111000100111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000111000101000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000111000101001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000111000101010" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000111000101111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000111000110000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000111000110001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000111000110010" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000111000110011" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000111000110100" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000111000110101" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000111000110110" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000111000110111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000111000111000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000111000111101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000111000111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111000111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111001000000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000111001000001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000111001000010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000111001000011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000111001000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111001000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111001000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111001000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111001001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111001001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111001001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111001001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111001001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111001001101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000111100100110" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000111100100111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000111100101001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000111100101010" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000111100111101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000111100111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111100111111" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0000111101000000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000111101000001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000111101000010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000111101000011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000111101000100" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0000111101000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111101000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111101000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111101001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111101001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111101001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111101001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000111101001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000000100101" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001000000100110" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001000000100111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001000000101000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0001000000101001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001000000101010" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001000000101011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001000000111101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001000000111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000000111111" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0001000001000000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0001000001000001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0001000001000010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0001000001000011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0001000001000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000001000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000001000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000001000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000001001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000001001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000001001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000001001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000001001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000100100100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0001000100100101" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001000100100110" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001000100100111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001000100101000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001000100101001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001000100101010" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001000100101011" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001000100111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000100111111" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0001000101000000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0001000101000001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0001000101000010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0001000101000011" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0001000101000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000101000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000101000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000101000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000101001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000101001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000101001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000101001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001000100100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001001000100101" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001001000100110" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001001000100111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001001000101000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001001000101001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001001000101010" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001001000101011" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001001000101100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001001000111110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001001000111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001001000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001001000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001001000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001001000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001001000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001001000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001001000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001001000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001001001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001001001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001001001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001100100100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001001100100101" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001001100100110" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001001100100111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001001100101000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001001100101001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001001100101010" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001001100101011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001001100101100" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001001100111111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001001101000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001101000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001101000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001101000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001101000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001101000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001101000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001101000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001101001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001101001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001010000100100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001010000100101" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001010000100110" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001010000100111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001010000101000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001010000101001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001010000101010" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001010000101011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001010000101100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001010000101101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001010001000001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001010001000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001010001000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001010001000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001010001000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001010001000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001010001000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001010100100100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001010100100101" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001010100100110" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001010100100111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001010100101000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001010100101001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001010100101010" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001010100101011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001010100101101" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001011000100101" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001011000100110" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001011000100111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001011000101000" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001011000101001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001011000101010" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001011000101011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001011000101110" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001011100100101" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001011100100110" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001011100100111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001011100101000" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001011100101001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001011100101010" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001011100101011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001011100101111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001100000100101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001100000100110" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001100000100111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001100000101000" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001100000101001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001100000101010" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001100000101011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0001100000101111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0001100000110000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001100000111011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001100000111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100000111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100000111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100000111111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001100001000000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001100100100110" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001100100100111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001100100101000" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001100100101001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001100100101010" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001100100110001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001100100111010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100100111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100100111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100100111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100100111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100100111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100101000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100101000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100101000010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001101000100110" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001101000100111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001101000101000" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001101000101001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001101000101010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001101000110010" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001101000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001101000111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0001101000111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101000111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101000111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101000111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101000111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101001000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101001000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101001000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101001000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101100100110" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001101100100111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001101100101000" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001101100101001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001101100110011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001101100110100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0001101100111000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001101100111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0001101100111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0001101100111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101100111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101100111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101100111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101100111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101101000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101101000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101101000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101101000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101101000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101110010001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001101110010010" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0001101110010011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0001101110010100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0001101110010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0001101110010110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0001101110010111" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0001101110011000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001110000100110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001110000100111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001110000101000" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001110000110101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001110000111000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110000111001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110000111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0001110000111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110000111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110000111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110000111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110000111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110001000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110001000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110001000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110001000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110001000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110001000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001110010001111" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0001110010010000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0001110010010001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001110010010010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001110010010011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0001110010010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001110010010101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001110010010110" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0001110010010111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001110010011000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001110010011001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0001110010011010" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0001110100100110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001110100100111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0001110100110110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0001110100110111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001110100111000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110100111001" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0001110100111010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001110100111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110100111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110100111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110100111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110100111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110101000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110101000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110101000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110101000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110101000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110101000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110110001101" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0001110110001110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0001110110001111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001110110010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001110110010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001110110010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001110110010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001110110010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001110110010101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001110110010110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001110110010111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001110110011000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001110110011001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001110110011010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001110110011011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0001110110011100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001111000100110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0001111000111000" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0001111000111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0001111000111010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111000111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111000111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111000111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111000111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111000111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111001000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111001000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111001000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111001000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111001000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111001000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111001000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001111010001100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0001111010001101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001111010001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111010001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111010010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111010010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111010010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111010010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111010010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111010010101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111010010110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111010010111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111010011000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111010011001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111010011010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111010011011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111010011100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0001111010011101" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0001111100110111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111100111000" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0001111100111001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111100111010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111100111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111100111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111100111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111100111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111100111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111101000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111101000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111101000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111101000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111101000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111101000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111101000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001111110001011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0001111110001100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001111110001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111110001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111110001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111110010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111110010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111110010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111110010011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0001111110010100" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0001111110010101" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0001111110010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001111110010111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001111110011000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111110011001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111110011010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111110011011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111110011100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001111110011101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001111110011110" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0010000000110110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010000000110111" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010000000111000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000000111001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000000111010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010000000111011" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010000000111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000000111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000000111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000000111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000001000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000001000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000001000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000001000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000001000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000001000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000001000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010000001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010000001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010000001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010000001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010000001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010000001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010000010001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0010000010001011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010000010001100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000010001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000010001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000010001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000010010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000010010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000010010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000010010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010000010010100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010000010010101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010000010010110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010000010010111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010000010011000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010000010011001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010000010011010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000010011011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000010011100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000010011101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000010011110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010000010011111" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0010000100110110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000100110111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000100111000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000100111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010000100111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010000100111011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010000100111100" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010000100111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000100111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000100111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000101000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000101000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000101000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000101000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000101000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000101000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000101000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010000101101011" => 
 	 	 	 	 color <= "111011";
 	 	 	when "0010000101101100" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010000101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010000101101110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010000101101111" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010000101110000" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010000110001001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0010000110001010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010000110001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000110001100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000110001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000110001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000110001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010000110010000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010000110010001" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010000110010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000110010011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010000110010100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010000110010101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010000110010110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010000110010111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010000110011000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010000110011001" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010000110011010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000110011011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000110011100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000110011101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000110011110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000110011111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0010001000110101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010001000110110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001000110111" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0010001000111000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010001000111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010001000111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010001000111011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010001000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010001000111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001000111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001000111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001001000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001001000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001001000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001001000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001001000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001001000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001001000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010001001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010001001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010001001101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010001010001000" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0010001010001001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010001010001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001010001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001010001100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001010001101" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010001010001110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001010001111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001010010000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001010010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010001010010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001010010011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001010010100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001010010101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001010010110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001010010111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001010011000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001010011001" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010001010011010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001010011011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001010011100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001010011101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001010011110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001010011111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001010100000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0010001100110101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010001100110110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001100110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010001100111000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010001100111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010001100111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010001100111011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010001100111100" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010001100111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001100111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001100111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001101000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001101000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001101000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001101000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001101000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001101000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001101000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010001101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010001101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010001101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010001110000111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0010001110001000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0010001110001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001110001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001110001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001110001100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010001110001101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001110001110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001110001111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001110010000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001110010001" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001110010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001110010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010001110010100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001110010101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001110010110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001110010111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001110011000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010001110011001" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010001110011010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001110011011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010001110011100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010001110011101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001110011110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001110011111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010001110100000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010001110100001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010010000110101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010010000110110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010000110111" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010010000111000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010010000111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010010000111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010010000111011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010010000111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010000111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010000111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010000111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010001000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010001000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010001000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010001000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010001000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010001000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010001000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010010001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010010001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010010001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010010001101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010010010000111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0010010010001000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010010010001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010010010001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010010010001011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010010010001100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010010001101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010010001110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010010001111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010010010000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010010010001" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010010010010" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010010010010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010010010100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010010010101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010010010110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010010010111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010010011000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010010011001" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010010010011010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010010011011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010010011100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010010011101" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010010010011110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010010010011111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010010010100000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010010010100001" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0010010100110110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010100110111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010100111000" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010010100111001" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010010100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010100111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010100111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010100111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010100111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010100111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010101000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010101000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010101000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010101000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010101000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010101000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010010101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010010101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010010101101100" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010010101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010010101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010010110000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010010110000111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0010010110001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010010110001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010010110001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010010110001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010010110001100" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010010110001101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010110001110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010110001111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010110010000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010110010001" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010110010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010110010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010110010100" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010010110010101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010110010110" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010010110010111" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010010110011000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010010110011001" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010110011010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010110011011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010110011100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010010110011101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010110011110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010010110011111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010010110100000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010010110100001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0010011000110110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010011000110111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011000111000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011000111001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011000111010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011000111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011000111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011000111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011000111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011000111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011001000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011001000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011001000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011001000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011001000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011001101010" => 
 	 	 	 	 color <= "100110";
 	 	 	when "0010011001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010011001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010011001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010011010000110" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0010011010000111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010011010001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010011010001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010011010001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010011010001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010011010001100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010011010001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010011010001110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010011010001111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010011010010000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010011010010001" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010011010010010" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010011010010011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010011010010100" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010011010010101" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010011010010110" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010011010010111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010011010011000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010011010011001" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010011010011010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010011010011011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010011010011100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010011010011101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010011010011110" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010011010011111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010011010100000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010011010100001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010011100110111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010011100111000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011100111001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011100111010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011100111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011100111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011100111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011100111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011100111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011101000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011101000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011101000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011101000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011101000100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010011101101010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010011101101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010011101101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010011101101101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010011101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010011101101111" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010011101110000" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010011110000110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0010011110000111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010011110001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010011110001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010011110001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010011110001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010011110001100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010011110001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010011110001110" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010011110001111" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010011110010000" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010011110010001" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010011110010010" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010011110010011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010011110010100" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010011110010101" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010011110010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010011110010111" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010011110011000" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010011110011001" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010011110011010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010011110011011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010011110011100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010011110011101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010011110011110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010011110011111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010011110100000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010011110100001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010011110100010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0010100000111000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010100000111001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100000111010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100000111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100000111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100000111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100000111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100000111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100001000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100001000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100001000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100001000011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010100001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010100001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010100001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010100001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010100001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010100001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010100001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010100010000110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0010100010000111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010100010001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010100010001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010100010001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100010001011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010100010001100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010100010001101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010100010001110" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010100010001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100010010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100010010001" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010100010010010" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010100010010011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010100010010100" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010100010010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100010010110" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010100010010111" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010100010011000" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010100010011001" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010100010011010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100010011011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100010011100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010100010011101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010100010011110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010100010011111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010100010100000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010100010100001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010100010100010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0010100100111010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010100100111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100100111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100100111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100100111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100100111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100101000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100101000001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010100101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010100101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010100101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010100101101110" => 
 	 	 	 	 color <= "100110";
 	 	 	when "0010100110000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010100110000110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010100110000111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010100110001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010100110001001" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010100110001010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010100110001011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010100110001100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010100110001101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010100110001110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010100110001111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010100110010000" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010100110010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100110010010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010100110010011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010100110010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010100110010101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010100110010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100110010111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100110011000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100110011001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010100110011010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100110011011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100110011100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100110011101" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010100110011110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100110011111" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010100110100000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010100110100001" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010100110100010" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0010101001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010101001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010101001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010101001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010101010000101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0010101010000110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010101010000111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010101010001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010101010001001" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010101010001010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101010001011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101010001100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101010001101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101010001110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101010001111" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010101010010000" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010101010010001" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010101010010010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010101010010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010101010010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010101010010101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010101010010110" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010101010010111" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010101010011000" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010101010011001" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101010011010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101010011011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101010011100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101010011101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101010011110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101010011111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010101010100000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010101010100001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010101010100010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0010101101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010101101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010101101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010101101101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010101101101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010101110000101" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0010101110000110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010101110000111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010101110001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010101110001001" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010101110001010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101110001011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101110001100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101110001101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101110001110" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010101110001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010101110010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010101110010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010101110010010" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010101110010011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010101110010100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010101110010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010101110010110" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010101110010111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010101110011000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101110011001" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101110011010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101110011011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101110011100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101110011101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101110011110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010101110011111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010101110100000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010101110100001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010101110100010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010110001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010110001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010110001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010110001101110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010110001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010110001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010110010000101" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0010110010000110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010110010000111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010110010001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010110010001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010110010001010" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010110010001011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010110010001100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010110010001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010110010001110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010110010001111" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010110010010000" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010110010010001" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010110010010010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010110010010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010110010010100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010110010010101" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010110010010110" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010110010010111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010110010011000" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010110010011001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010110010011010" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010110010011011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010110010011100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010110010011101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010110010011110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010110010011111" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010110010100000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010110010100001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010110101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010110101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010110101101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010110101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010110101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010110101101111" => 
 	 	 	 	 color <= "010001";
 	 	 	when "0010110101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010110110000101" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0010110110000110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010110110000111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010110110001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010110110001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010110110001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010110110001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010110110001100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010110110001101" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010110110001110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010110110001111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010110110010000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010110110010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010110110010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010110110010011" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010110110010100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010110110010101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010110110010110" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010110110010111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010110110011000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010110110011001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010110110011010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010110110011011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010110110011100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010110110011101" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010110110011110" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010110110011111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010110110100000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010110110100001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0010111001101010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010111001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010111001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010111001101101" => 
 	 	 	 	 color <= "111011";
 	 	 	when "0010111001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010111010000101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0010111010000110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010111010000111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111010001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111010001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111010001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111010001011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010111010001100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111010001101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111010001110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111010001111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111010010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010111010010001" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010111010010010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111010010011" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010111010010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010111010010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010111010010110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111010010111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111010011000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111010011001" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010111010011010" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010111010011011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111010011100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111010011101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111010011110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111010011111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111010100000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111010100001" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0010111101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010111101101100" => 
 	 	 	 	 color <= "101011";
 	 	 	when "0010111101101101" => 
 	 	 	 	 color <= "101011";
 	 	 	when "0010111101101110" => 
 	 	 	 	 color <= "101011";
 	 	 	when "0010111101101111" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010111101110000" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010111110000110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0010111110000111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111110001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111110001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111110001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111110001011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010111110001100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111110001101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111110001110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111110001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010111110010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111110010001" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0010111110010010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111110010011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111110010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010111110010101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010111110010110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111110010111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111110011000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111110011001" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111110011010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0010111110011011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010111110011100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111110011101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111110011110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111110011111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010111110100000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010111110100001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0011000001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011000001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011000001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011000001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011000001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011000001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011000001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011000010000110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011000010000111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0011000010001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000010001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000010001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000010001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000010001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011000010001101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000010001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011000010001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000010010000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0011000010010001" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000010010010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000010010011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000010010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011000010010101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000010010110" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000010010111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000010011000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000010011001" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000010011010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000010011011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000010011100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0011000010011101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000010011110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000010011111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000010100000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011000101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011000101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011000101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011000101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011000101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011000110000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0011000110000111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011000110001000" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0011000110001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000110001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000110001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000110001100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0011000110001101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0011000110001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000110001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000110010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011000110010001" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000110010010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000110010011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000110010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011000110010101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000110010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011000110010111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000110011000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000110011001" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000110011010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000110011011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011000110011100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0011000110011101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000110011110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000110011111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0011000110100000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0011001001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011001001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011001001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011001001101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011001001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011001010000111" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0011001010001000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011001010001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001010001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001010001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001010001100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001010001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001010001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001010001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001010010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011001010010001" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011001010010010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011001010010011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011001010010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011001010010101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001010010110" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0011001010010111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011001010011000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011001010011001" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011001010011010" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0011001010011011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0011001010011100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001010011101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001010011110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001010011111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011001101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011001101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011001101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011001101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011001101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011001110001000" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0011001110001001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011001110001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001110001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001110001100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001110001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001110001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001110001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001110010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001110010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011001110010010" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011001110010011" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0011001110010100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0011001110010101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001110010110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001110010111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011001110011000" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0011001110011001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0011001110011010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001110011011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001110011100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001110011101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011001110011110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011001110011111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0011010001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011010001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011010001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011010001101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011010001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011010010001001" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0011010010001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011010010001011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0011010010001100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010010101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010010110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010010111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010011000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010011001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010011010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010011011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010011100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010010011101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011010010011110" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0011010101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011010101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011010101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011010101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011010101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011010110001010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0011010110001011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011010110001100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011010110001101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0011010110001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010110001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010110010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010110010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010110010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010110010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010110010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010110010101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010110010110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010110010111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010110011000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010110011001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010110011010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010110011011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0011010110011100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011010110011101" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0011011001101010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011011001101011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011011001101101" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011011001101110" => 
 	 	 	 	 color <= "010001";
 	 	 	when "0011011001110000" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011011010001100" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0011011010001101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011011010001110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011011010001111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0011011010010000" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0011011010010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011011010010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011011010010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011011010010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011011010010101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011011010010110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011011010010111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011011010011000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011011010011001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0011011010011010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011011010011011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011011010011100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0011011101101010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011011101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011011101101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011011101101101" => 
 	 	 	 	 color <= "101111";
 	 	 	when "0011011101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011011110001110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0011011110001111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011011110010000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011011110010001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011011110010010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011011110010011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011011110010100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0011011110010101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0011011110010110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011011110010111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011011110011000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011011110011001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0011011110011010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0011100001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011100001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011100001101100" => 
 	 	 	 	 color <= "111011";
 	 	 	when "0011100001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011100001101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011100001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011100010010001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0011100010010010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0011100010010011" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0011100010010100" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0011100010010101" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0011100010010110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0011100010010111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0011100101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011100101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011100101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011100101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011100101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011101000111101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0011101000111110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0011101000111111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0011101001010100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0011101001010101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0011101001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011101001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011101001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011101001101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011101001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011101100111011" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0011101100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011101100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011101100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011101100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011101101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011101101000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011101101010001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0011101101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011101101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011101101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011101101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011101101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011101101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011101101011000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0011101101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011101101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011101101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011101101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011101101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011110000111010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011110000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110001000011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0011110001010000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0011110001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110001011001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0011110001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011110001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011110001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011110001101110" => 
 	 	 	 	 color <= "011010";
 	 	 	when "0011110001101111" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011110001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011110100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011110101000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0011110101001111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0011110101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011110101011010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0011110101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011110101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011110101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011110101101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011110101101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011110101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011111000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111001000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0011111001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111001011011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0011111001101010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011111001101011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011111001101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011111001101111" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011111001110000" => 
 	 	 	 	 color <= "010001";
 	 	 	when "0011111100111000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0011111100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011111101001110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0011111101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0011111101101010" => 
 	 	 	 	 color <= "011010";
 	 	 	when "0011111101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011111101101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011111101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0011111101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100000000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000001001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000001001010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0100000001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001011100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0100000001100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000001100011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100000001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100000001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100000001101100" => 
 	 	 	 	 color <= "100110";
 	 	 	when "0100000001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100000001101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0100000001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100000100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000101001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000101001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000101001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100000101001100" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0100000101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000101010011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100000101010100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100000101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000101011100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0100000101011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100000101100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000101100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000101100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000101100011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100000101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100000101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0100000101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100000101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0100000101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100001000110111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100001000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001001001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001001001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001001001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001001001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001001001101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0100001001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001001010010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100001001010011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100001001010100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100001001010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100001001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001001011100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100001001011101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100001001011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100001001100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001001100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001001100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001001100011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001001100100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100001001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100001001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0100001001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100001001101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0100001001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100001100110111" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0100001100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001101001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001101001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001101001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001101001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001101001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100001101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001101010011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100001101010101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100001101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001101011100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100001101011101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100001101011111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0100001101100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001101100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001101100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001101100011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001101100100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100001101100101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100001101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100001101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0100001101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100001101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0100001101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100010000110111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100010000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010000111110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100010000111111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100010001000000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100010001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010001001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010001001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010001001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010001001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010001001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001011101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0100010001011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100010001100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001100011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001100100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010001100101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100010001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100010001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0100010001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100010001101110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0100010001101111" => 
 	 	 	 	 color <= "011010";
 	 	 	when "0100010001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100010100111000" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0100010100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010100111101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100010100111110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100010100111111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100010101000000" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0100010101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010101001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010101001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010101001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010101001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010101001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100010101001110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0100010101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101010011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100010101010100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100010101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101100011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101100100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100010101100101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100010101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100010101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0100010101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100010101101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100010101101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100010101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100011000111001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100011000111010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0100011000111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100011000111100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100011000111101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100011000111110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100011000111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100011001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011001001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011001001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011001001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011001001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011001001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011001001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011001001111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0100011001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011001010001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0100011001010010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100011001010011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100011001010100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100011001010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100011001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011001011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011001100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011001100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011001100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011001100011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011001100100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011001100101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100011100111011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100011100111100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100011100111101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100011100111111" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0100011101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011101000111" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0100011101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011101001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011101001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011101001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011101001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011101001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011101001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011101001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100011101010000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0100011101010001" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0100011101010010" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100011101010011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100011101010100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100011101010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100011101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011101100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011101100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011101100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011101100011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100011101100100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100011101100101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100100000111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100100001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100001000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100100001001000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100100001001001" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0100100001001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100001001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100001001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100001001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100001001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100001001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100001010000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100100001010001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100100001010110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100100001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100001011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100001100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100001100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100001100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100001100011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100001100100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0100100001100101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100100100110111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100100100111000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100100100111001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100100101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100101000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100100101000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100100101001000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100100101001010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100100101001011" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0100100101001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100101001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100101001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100101001111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100100101010000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100100101010001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100100101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100101100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100101100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100101100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100101100011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100100101100100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100100101100101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100101000110101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100101000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101000111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100101000111111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100101001000000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100101001000001" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0100101001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101001000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100101001000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100101001000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100101001001100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100101001001101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100101001001110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100101001001111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100101001010000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100101001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101001011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101001100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101001100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101001100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101001100011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0100101001100100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100101001100101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100101001101011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0100101001101100" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0100101001101101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0100101001101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0100101001101111" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0100101001110000" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0100101100110100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100101100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100101101000011" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0100101101000100" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0100101101000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100101101000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100101101000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100101101001110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100101101001111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0100101101010000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0100101101010001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0100101101010010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100101101010011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100101101010100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100101101010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100101101010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100101101010111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100101101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101101100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101101100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100101101100010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0100101101100011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100101101100100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100101101101010" => 
 	 	 	 	 color <= "101111";
 	 	 	when "0100101101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100101101101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100101101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100101101101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100101101101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100101101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100110000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110001001000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100110001001101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100110001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110001100000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100110001100001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100110001100010" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100110001100011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100110001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100110001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0100110001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100110001101110" => 
 	 	 	 	 color <= "100110";
 	 	 	when "0100110100110011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100110100110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110101001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100110101001010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0100110101001011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100110101001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100110101011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0100110101100000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100110101100001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100110101100010" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0100110101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100110101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0100110101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100110101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0100111000110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111001001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111001001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111001100000" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0100111001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100111001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0100111001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100111001101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0100111100110010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100111100110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111100110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100111101001001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0100111101001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0100111101100001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0100111101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100111101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0100111101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100111101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101000000110010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101000000110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000001001001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000001100001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0101000001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000001110111" => 
 	 	 	 	 color <= "011010";
 	 	 	when "0101000001111000" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101000001111001" => 
 	 	 	 	 color <= "011010";
 	 	 	when "0101000001111100" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101000001111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101000100110010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0101000100110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000100110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000100111001" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0101000100111010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101000100111011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101000100111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101000100111101" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0101000100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000101001001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101000101100001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0101000101100010" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101000101101010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101000101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000101101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000101101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000101101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000101110110" => 
 	 	 	 	 color <= "011010";
 	 	 	when "0101000101110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000101111000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000101111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000101111010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101000101111100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000101111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101001000110010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001000110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001000111001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101001000111010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101001000111011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101001000111101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101001000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001001001001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001001111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101001001010000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101001001010001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101001001010010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101001001010011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101001001010100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0101001001010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0101001001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001001100001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101001001100010" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101001001101010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101001001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101001001101100" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101001001101101" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101001001101110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101001001101111" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101001001110000" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101001001110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101001001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101001001111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101001001111010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101001001111100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101001001111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101001100110010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001100110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001100110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001100111010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101001100111100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101001100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101001101001001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101010001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0101001101010010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0101001101010011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101001101010100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101001101010101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101001101010110" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0101001101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101001101100000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101001101100001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101001101100010" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101001101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101001101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101001101101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101001101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101001101101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101001101101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101001101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101001101110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101001101110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101001101111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101001101111010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101001101111100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101001101111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101010000110010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0101010000110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010001000110" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0101010001000111" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0101010001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010001001001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0101010001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010001011100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101010001011101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101010001011110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101010001011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101010001100000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101010001100001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101010001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101010001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101010001101101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101010001110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101010001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101010001111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101010001111010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101010001111100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101010001111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101010100110010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101010100110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010100110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101010101000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101010101001000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101010101001001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0101010101001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101010101011100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101010101011101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101010101101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101010101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101010101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101010101110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101010101110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101010101111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101010101111010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101010101111100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101010101111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101011000110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011001001000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101011001001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011001011100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0101011001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101011001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101011001101111" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101011001110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101011001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101011001111001" => 
 	 	 	 	 color <= "111011";
 	 	 	when "0101011001111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101011001111011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101011001111100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101011001111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101011100110011" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0101011100110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101011101001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101011101101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101011101101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101011101110000" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101011101110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101011101110111" => 
 	 	 	 	 color <= "111011";
 	 	 	when "0101011101111010" => 
 	 	 	 	 color <= "111011";
 	 	 	when "0101011101111011" => 
 	 	 	 	 color <= "111011";
 	 	 	when "0101011101111100" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101100000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100001001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100001001100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0101100001001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100001011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0101100001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101100001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101100001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101100001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101100001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101100001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101100001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101100001110110" => 
 	 	 	 	 color <= "011010";
 	 	 	when "0101100001110111" => 
 	 	 	 	 color <= "101111";
 	 	 	when "0101100100110101" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0101100100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100100111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101100101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100101001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100101001010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101100101001101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101100101001110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0101100101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101100101011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0101100101011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101100101101010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101100101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101100101101100" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101100101101101" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101100101101110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101100101101111" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101100101110000" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101100101110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101100101110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101101000110110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101000110111" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0101101000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101000111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101101000111110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101000111111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101001000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101101001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101001001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101001001010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101001001111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101101001010000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0101101001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101001011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0101101001011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101101001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101101001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101101001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101101001101101" => 
 	 	 	 	 color <= "101111";
 	 	 	when "0101101001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101101001110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101101001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101101100001101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101100001110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101101100001111" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0101101100010000" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0101101100010001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101101100010010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101100111000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101100111001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101100111010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101100111011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101100111100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101100111101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101100111110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101100111111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101101000001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101101101001001" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0101101101001010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101101001011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101101101010000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101101101010001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0101101101010010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0101101101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101101101011110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101101101011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101101101101010" => 
 	 	 	 	 color <= "111011";
 	 	 	when "0101101101101011" => 
 	 	 	 	 color <= "111011";
 	 	 	when "0101101101101100" => 
 	 	 	 	 color <= "111011";
 	 	 	when "0101101101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101101101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101101101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101101101110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101101101110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101101101111000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101101101111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101101101111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101101101111011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101101101111100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101101101111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101110000001010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101110000001011" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0101110000001100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101110000001101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101110000001110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101110000001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0101110000010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0101110000010001" => 
 	 	 	 	 color <= "111101";
 	 	 	when "0101110000010010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101110000010011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101110000010100" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0101110000010101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101110000111001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101110000111010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101110000111011" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0101110000111100" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0101110000111101" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0101110000111110" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0101110000111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101110001000000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101110001000001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101110001000010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101110001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110001001001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101110001001010" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0101110001001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110001011101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101110001011110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101110001011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101110001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101110001101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101110001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101110001110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101110001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101110001111000" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101110001111001" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101110001111010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101110001111011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101110001111100" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101110001111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101110100001001" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0101110100001010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101110100001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0101110100001100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101110100001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0101110100001110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101110100001111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101110100010000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101110100010001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101110100010010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101110100010011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101110100010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0101110100010101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101110100010110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101110100110100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101110100110101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101110100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101110101001000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101110101001001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101110101011101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101110101011110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0101110101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101110101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101110101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101110101110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101110101110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101111000000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101111000001000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101111000001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0101111000001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0101111000001011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101111000001100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0101111000001101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101111000001110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101111000001111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101111000010000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101111000010001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101111000010010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101111000010011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101111000010100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101111000010101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0101111000010110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0101111000010111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101111000011000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101111000110010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101111000110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111001000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101111001000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101111001001000" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0101111001001001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101111001101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101111001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101111001110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0101111001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101111100000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101111100000111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101111100001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0101111100001001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101111100001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101111100001011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101111100001100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101111100001101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101111100001110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101111100001111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101111100010000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101111100010001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101111100010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0101111100010011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101111100010100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101111100010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0101111100010110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101111100010111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0101111100011000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0101111100011001" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0101111100110001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101111100110010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111100110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111100110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101111101000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101111101001000" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0101111101001001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0101111101011110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0101111101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101111101101110" => 
 	 	 	 	 color <= "011010";
 	 	 	when "0101111101101111" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0101111101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101111101110110" => 
 	 	 	 	 color <= "010001";
 	 	 	when "0101111101110111" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110000000000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110000000000110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110000000000111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000000001000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110000000001001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000000001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000000001011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000000001100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000000001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110000000001110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000000001111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000000010000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000000010001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000000010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110000000010011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000000010100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000000010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000000010110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000000010111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110000000011000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000000011001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110000000011010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110000000110001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000000110010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000000110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000001001000" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0110000001001001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000001011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110000001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000001111000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000001111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000001111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000001111011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000001111100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000001111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110000100000101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000100000110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110000100000111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110000100001000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000100001001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000100001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000100001011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000100001100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000100001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110000100001110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000100001111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000100010000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000100010001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110000100010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110000100010011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000100010100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000100010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000100010110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000100010111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000100011000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110000100011001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110000100011010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110000100110001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000100110010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000100110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000100110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000101001000" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0110000101001001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110000101011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110000101011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110000101101010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110000101101011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110000101101100" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110000101101101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110000101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110000101101111" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110000101110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110000101110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000101111000" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110000101111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000101111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000101111011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110000101111100" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110000101111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110001000000100" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0110001000000101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110001000000110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110001000000111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110001000001000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110001000001001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001000001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001000001011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001000001100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001000001101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110001000001110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110001000001111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001000010000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001000010001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110001000010010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110001000010011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001000010100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001000010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001000010110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001000010111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110001000011000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110001000011001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110001000011010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110001000011011" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0110001000110001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001000110010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001000110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001001001001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0110001001001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001001011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110001001011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110001001110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110001001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110001001111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110001001111010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110001100000100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001100000101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110001100000110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110001100000111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001100001000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110001100001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110001100001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001100001011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001100001100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001100001101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001100001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110001100001111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001100010000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001100010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110001100010010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001100010011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001100010100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001100010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001100010110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110001100010111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110001100011000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001100011001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001100011010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110001100011011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110001100110001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001100110010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001100110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001100110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110001101001001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110001101001010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0110001101001011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0110001101001100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0110001101001101" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0110001101001110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110001101001111" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0110001101010000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0110001101010001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0110001101010010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0110001101010011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110001101010100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110001101010101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110001101010110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110001101010111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110001101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110001101011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110001101011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110001101110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110001101110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110001101111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110001101111010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110010000000011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010000000100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110010000000101" => 
 	 	 	 	 color <= "111101";
 	 	 	when "0110010000000110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010000000111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010000001000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010000001001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110010000001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110010000001011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110010000001100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010000001101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010000001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110010000001111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010000010000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010000010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110010000010010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010000010011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010000010100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110010000010101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110010000010110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110010000010111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010000011000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010000011001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010000011010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110010000011011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110010000011100" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0110010000110010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010000110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010000111000" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0110010000111001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110010000111010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010000111011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010000111100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010000111101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010000111110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010000111111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010001001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110010001001010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010001001100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110010001001101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110010001001110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110010001001111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110010001010000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110010001010001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110010001010010" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110010001010011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110010001010100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110010001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110010001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110010001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110010001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110010001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110010001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110010001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110010001011110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0110010001011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110010001110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110010001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110010001111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110010001111010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110010100000011" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0110010100000100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110010100000101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110010100000110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010100000111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010100001000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010100001001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010100001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010100001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110010100001100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110010100001101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010100001110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110010100001111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110010100010000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110010100010001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110010100010010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010100010011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110010100010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110010100010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010100010110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010100010111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010100011000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010100011001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010100011010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110010100011011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110010100011100" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0110010100110011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010100110100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010100110101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010100110110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010100110111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010100111000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010100111001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010100111010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010100111011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010100111100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010100111101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110010101001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110010101001010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110010101010111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110010101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110010101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110010101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110010101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110010101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110010101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110010101011110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110010101011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110010101110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110010101110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110010101111000" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110010101111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110010101111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110010101111011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110010101111100" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110011000000011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000000100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110011000000101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000000110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000000111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000001000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000001001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000001011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000001100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110011000001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110011000001110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110011000010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110011000010001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110011000010011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110011000010100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000010110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000010111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000011000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000011001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000011010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000011011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110011000011100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011000110101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110011000110110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110011000110111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110011000111000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110011000111111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110011001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011001001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110011001001010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110011001010111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0110011001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110011001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110011001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110011001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110011001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110011001011101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110011001011110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110011001011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110011001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011001110110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110011001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011001111000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011001111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011001111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011001111011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011001111100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011001111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110011100000011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100000100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011100000101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110011100000110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100000111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100001000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100001001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100001011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100001100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100001101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110011100001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110011100001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110011100010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110011100010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110011100010010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110011100010011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100010100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100010110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100010111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100011000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100011001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100011010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100011011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011100011100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110011100111000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110011100111001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110011100111010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110011100111011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110011100111100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110011100111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110011100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110011101001001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110011101001010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110011101010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110011101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110011101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110011101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110011101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110011101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110011101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110011101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110011101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110011101011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110011101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011101101100" => 
 	 	 	 	 color <= "100110";
 	 	 	when "0110011101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011101101110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110011101101111" => 
 	 	 	 	 color <= "100110";
 	 	 	when "0110011101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110011101110111" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110011101111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110011101111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110011101111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110011101111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110011101111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110011101111101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0110100000000011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100000000100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100000000101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100000000110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000000111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000001100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000001111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100000010000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100000010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000010101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000010110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000010111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000011000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000011001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100000011010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100000011011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100000011100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110100000110011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110100000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100001001001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110100001001010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110100001010010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0110100001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110100001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100001101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110100001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100001110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110100001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100001111000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100001111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100001111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100001111011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100001111100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100001111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110100100000011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100000100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100100000101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110100100000110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100000111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100001000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100001001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100001011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100001100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100001101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100100001111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100100010000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100100010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110100100010010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110100100010011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100010100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100010110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100010111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100011000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100011001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100011010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110100100011011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100100011100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110100100110001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110100100110010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100100110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100100110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110100101001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110100101001001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110100101001010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110100101010000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0110100101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110100101011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110100101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110100101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110100101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100101110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110100101110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100101111000" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110100101111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100101111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110100101111011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110100101111100" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110101000000011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000000100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110101000000101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000000110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000000111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000001000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000001001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000001011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000001100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110101000001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110101000001110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110101000001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110101000010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110101000010001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110101000010011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110101000010100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000010110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000010111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000011000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000011001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000011010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000011011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110101000011100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101000110001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101000110010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101000110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101001001000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110101001001001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110101001001110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110101001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101001011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110101001100000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110101001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110101001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110101001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110101001101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110101001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110101001110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110101001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110101001111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110101001111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110101100000011" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0110101100000100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110101100000101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101100000110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101100000111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101100001000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101100001001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101100001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101100001011" => 
 	 	 	 	 color <= "111101";
 	 	 	when "0110101100001100" => 
 	 	 	 	 color <= "111101";
 	 	 	when "0110101100001101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101100001110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110101100001111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110101100010000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110101100010001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110101100010010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101100010011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110101100010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110101100010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101100010110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101100010111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101100011000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101100011001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101100011010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110101100011011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110101100011100" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0110101100110000" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0110101100110001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101100110010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101100110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101100110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110101101000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110101101001000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110101101001001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110101101001101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110101101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110101101011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110101101100000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110101101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110101101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110101101101100" => 
 	 	 	 	 color <= "011010";
 	 	 	when "0110101101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110101101101110" => 
 	 	 	 	 color <= "101111";
 	 	 	when "0110101101101111" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110101101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110101101110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110101101110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110101101111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110101101111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110101101111011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110110000000011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110110000000100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110110000000101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110110000000110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110000000111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110000001000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110000001001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110110000001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110110000001011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110110000001100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110000001101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110000001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110110000001111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110000010000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110000010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110110000010010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110000010011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110000010100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110110000010101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110110000010110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110110000010111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110000011000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110000011001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110000011010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110110000011011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110110000011100" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0110110000110000" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0110110000110001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110000110010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110000110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110001000101" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0110110001000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110110001000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110110001001000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110110001001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110001011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110110001011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110110001100000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110110001101010" => 
 	 	 	 	 color <= "100110";
 	 	 	when "0110110001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110110001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110110001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110110001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110110001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110110001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110110001110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110110001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110110001111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110110001111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110110001111011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110110001111100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110110100000100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110100000101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110110100000110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110110100000111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110100001000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110110100001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110110100001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110100001011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110100001100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110100001101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110100001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110110100001111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110100010000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110100010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110110100010010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110100010011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110100010100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110100010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110100010110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110110100010111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110110100011000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110100011001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110100011010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110110100011011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110110100110000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110110100110001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110100110010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110100110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110100110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110110101000011" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0110110101000100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110110101000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110110101000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110110101000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110110101001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110110101011100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110110101011101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0110110101011110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110110101011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110110101100000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110110101101010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110110101101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110110101101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110110101101101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110110101101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110110101101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110110101110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110110101110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110110101111000" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110110101111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110110101111010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0110110101111100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110110101111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110111000000100" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0110111000000101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110111000000110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110111000000111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110111000001000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110111000001001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111000001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111000001011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111000001100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111000001101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110111000001110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110111000001111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111000010000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111000010001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110111000010010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110111000010011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111000010100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111000010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111000010110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111000010111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110111000011000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110111000011001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110111000011010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110111000011011" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0110111000110001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110111000110010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111000110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111001000001" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0110111001000010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110111001000011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110111001000100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110111001000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110111001000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110111001001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111001011100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110111001011101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110111001011110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0110111001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110111001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110111001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110111001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110111001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110111001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110111001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110111001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110111001111000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110111001111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110111001111010" => 
 	 	 	 	 color <= "010001";
 	 	 	when "0110111001111100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110111001111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110111100000101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111100000110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110111100000111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110111100001000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111100001001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111100001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111100001011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111100001100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111100001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110111100001110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111100001111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111100010000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111100010001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110111100010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110111100010011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111100010100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111100010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111100010110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111100010111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111100011000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0110111100011001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110111100011010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0110111100110010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0110111100110011" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0110111100110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111100111100" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0110111100111101" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0110111100111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110111100111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110111101000000" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0110111101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110111101001000" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0110111101001001" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0110111101001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111101001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111101001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111101001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111101010100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0110111101010101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0110111101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0110111101011100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0110111101101111" => 
 	 	 	 	 color <= "010001";
 	 	 	when "0110111101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110111101110110" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0110111101110111" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0111000000000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111000000000110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111000000000111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111000000001000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111000000001001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000000001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000000001011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000000001100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000000001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111000000001110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000000001111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000000010000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000000010001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000000010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111000000010011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000000010100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000000010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000000010110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000000010111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000000011000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111000000011001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111000000011010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111000000110100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111000000110101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111000000110110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111000000110111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111000000111000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111000000111001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111000000111010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111000000111011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111000000111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0111000000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000001001001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000001001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000001001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000001001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000001001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000001010001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111000001010010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0111000001010011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111000001010100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111000001010101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111000001010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111000001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000001011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111000001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111000001110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111000001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111000100000110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0111000100000111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111000100001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111000100001001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111000100001010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000100001011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000100001100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111000100001101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111000100001110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000100001111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000100010000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000100010001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000100010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111000100010011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111000100010100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000100010101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111000100010110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111000100010111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111000100011000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111000100011001" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0111000100110111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111000100111000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111000100111001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111000100111010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0111000100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111000101001001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101001111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0111000101010000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0111000101010001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0111000101010010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111000101010011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111000101010100" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0111000101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111000101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111000101110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111000101110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111001000000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111001000001000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111001000001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111001000001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111001000001011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111001000001100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111001000001101" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111001000001110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111001000001111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111001000010000" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111001000010001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111001000010010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111001000010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111001000010100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111001000010101" => 
 	 	 	 	 color <= "111101";
 	 	 	when "0111001000010110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111001000010111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111001000011000" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0111001000110111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111001000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001001001001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001001100000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111001001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111001001110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111001001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111001001111000" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111001001111001" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111001001111010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111001001111011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111001001111100" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111001001111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0111001100001001" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111001100001010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111001100001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111001100001100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111001100001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111001100001110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111001100001111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111001100010000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111001100010001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111001100010010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111001100010011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111001100010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111001100010101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111001100010110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111001100010111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111001100110101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111001100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111001101001001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111001101100001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111001101101010" => 
 	 	 	 	 color <= "101111";
 	 	 	when "0111001101101011" => 
 	 	 	 	 color <= "101111";
 	 	 	when "0111001101101100" => 
 	 	 	 	 color <= "101111";
 	 	 	when "0111001101101101" => 
 	 	 	 	 color <= "101111";
 	 	 	when "0111001101101110" => 
 	 	 	 	 color <= "101111";
 	 	 	when "0111001101101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111001101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111001101110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111001101110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111001101111000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111001101111001" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111001101111010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111001101111011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111001101111100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111001101111101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0111010000001010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111010000001011" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0111010000001100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111010000001101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111010000001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111010000001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111010000010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111010000010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0111010000010010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111010000010011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111010000010100" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0111010000010101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111010000110100" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0111010000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010001001001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0111010001001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010001100000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111010001100001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111010001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111010001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111010001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111010001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111010001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111010001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111010001110000" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111010001110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111010001110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111010100001101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111010100001110" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0111010100001111" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0111010100010000" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0111010100010001" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0111010100010010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111010100110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111010101001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0111010101001010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111010101100000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111010101100001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111010101101010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111010101101011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0111010101110110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111010101110111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111011000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011001000111" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0111011001001000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111011001001001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111011001001010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0111011001001011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011001100001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111011001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111011001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111011001110110" => 
 	 	 	 	 color <= "100110";
 	 	 	when "0111011001110111" => 
 	 	 	 	 color <= "111011";
 	 	 	when "0111011100110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111011101000100" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0111011101000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0111011101000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111011101000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111011101001000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111011101001001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111011101001100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101001101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111011101100010" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111011101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111011101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111100000110100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100000110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100001000001" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0111100001000010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111100001000011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111100001000100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111100001000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111100001000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111100001000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111100001001101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0111100001001110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111100001001111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111100001010000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111100001010001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111100001010010" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0111100001010011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111100001010100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111100001010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111100001010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111100001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100001011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100001100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100001100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100001100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111100001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111100001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111100001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111100001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111100001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111100001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111100100110100" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0111100100110101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111100100111100" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0111100100111101" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0111100100111110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111100100111111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111100101000000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111100101000001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111100101000010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111100101000011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111100101000100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111100101000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111100101001111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111100101010000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111100101010001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111100101010010" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111100101010011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111100101010100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0111100101010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111100101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100101100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100101100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100101100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111100101100011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111100101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111100101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111100101101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111100101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111100101101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111100101101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111100101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111101000110101" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0111101000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111101000110111" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0111101000111000" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0111101000111001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101000111010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101000111011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101000111100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101000111101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101000111110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101000111111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101001000000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101001000001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101001001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0111101001001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111101001001011" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0111101001001100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101001010010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0111101001010011" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0111101001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101001011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101001100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101001100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101001100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101001100011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111101001100100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111101001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111101001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111101100110110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101100110111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101100111000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101100111001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101100111010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101100111011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101100111100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101101000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111101101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111101101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111101101001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111101101001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111101101001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111101101001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111101101001101" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0111101101010000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111101101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111101101100011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111101101100100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111101101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111101101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111110000110111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111110000111000" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0111110000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110000111010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0111110001000100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111110001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110001001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110001001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110001001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110001001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110001001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110001001110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0111110001001111" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0111110001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110001100011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111110001100100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111110001101010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111110001101011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0111110100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110100111100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111110101000010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111110101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110101001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110101001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110101001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110101001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111110101001101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0111110101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101011010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111110101011011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111110101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111110101100011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111110101100100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111110101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111110101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111111000110110" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0111111000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111001000000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111111001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111001001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111001001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111001001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111001001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111001001101" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0111111001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001011000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111111001011001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0111111001011010" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111111001011011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111111001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111001100011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0111111001100100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111111001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111111001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0111111100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111100111101" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0111111100111110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111111100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111101001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111101001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111101001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111101001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0111111101001101" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0111111101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111101010101" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0111111101010110" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0111111101010111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111111101011000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111111101011001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111111101011010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0111111101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111101100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111101100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111101100010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0111111101100011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111111101100100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0111111101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0111111101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1000000000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000001001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000001001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000001001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000001001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000001001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000001001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000001010101" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1000000001010110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000000001010111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000000001011000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000000001011001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000000001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000001011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000001100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000001100001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000001100010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000000001100011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000000001100100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000000001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000000001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000000001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000000001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000000001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000000001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000000001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000000100110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000101001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000101001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000101001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000101001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000000101001101" => 
 	 	 	 	 color <= "100100";
 	 	 	when "1000000101001110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000000101100001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1000000101100010" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000000101100011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000000101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000000101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000000101101100" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1000000101101101" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1000000101101110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1000000101101111" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1000000101110000" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1000001000110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001001000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001001001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001001001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001001001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001001001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001001001100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000001001001101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000001001001110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1000001001001111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001100000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001001100001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1000001001100010" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000001001100011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000001001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000001001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1000001010001100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000001010001101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000001010001110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1000001100110110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1000001100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001101000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001101000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001101000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001101000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001101001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001101001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000001101001010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000001101001011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000001101001100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000001101001101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000001101001110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000001101001111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000001101010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001101011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001101011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001101011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000001101100000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1000001101100001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000001101100010" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000001101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000001101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1000001110001011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1000001110001100" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1000001110001101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000001110001110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000001110001111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000010000110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010001000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010001000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010001000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010001000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010001000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010001000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1000010001001000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000010001001001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000010001001010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000010001001011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000010001001100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000010001010000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010001010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010001010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010001011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010001011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010001011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010001011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010001011111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1000010001100000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000010001100001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000010001101010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1000010001101011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1000010010001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000010010001100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000010010001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000010010001110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000010010001111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000010010010000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000010010010001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000010100110111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000010101000011" => 
 	 	 	 	 color <= "100101";
 	 	 	when "1000010101000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1000010101000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000010101000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000010101000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000010101001000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000010101001001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000010101001010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000010101010001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010101010010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010101010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010101010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010101010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010101010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010101010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010101011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010101011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010101011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010101011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010101011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000010101011101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000010101011110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000010101011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000010101100000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000010101101010" => 
 	 	 	 	 color <= "011010";
 	 	 	when "1000010101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000010101101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000010101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000010101101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000010101101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000010101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000010110001010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "1000010110001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000010110001100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000010110001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000010110001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000010110001111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000010110010000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000010110010001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000011000110111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000011000111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011001000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1000011001000010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000011001000011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000011001000100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000011001000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000011001000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000011001000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000011001010010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000011001010011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000011001010100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000011001010101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000011001010110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000011001010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000011001011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000011001011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000011001011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "1000011001011011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000011001011100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1000011001011101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000011001011110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000011001011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000011001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000011001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000011001101100" => 
 	 	 	 	 color <= "100110";
 	 	 	when "1000011001101101" => 
 	 	 	 	 color <= "100110";
 	 	 	when "1000011001101110" => 
 	 	 	 	 color <= "100110";
 	 	 	when "1000011001101111" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1000011001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000011010001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011010001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011010001100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "1000011010001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000011010001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000011010001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000011010010000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000011010010001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000011010010010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000011100111000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011101000010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000011101000011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000011101010011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000011101010100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1000011101010101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1000011101010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000011101010111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000011101011000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1000011101011001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1000011101011010" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000011101011011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000011101011100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000011101011101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000011101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000011101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1000011101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000011110001001" => 
 	 	 	 	 color <= "100001";
 	 	 	when "1000011110001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011110001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011110001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011110001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000011110001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000011110001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000011110010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000011110010001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000011110010010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000011110010011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000100000111000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000100000111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100001000010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000100001010110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000100001010111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000100001011000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000100001011001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000100001011010" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000100001011011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1000100001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000100001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1000100001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000100010001000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000100010001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100010001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100010001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100010001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100010001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100010001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100010001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000100010010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000100010010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000100010010010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000100010010011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000100010010100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1000100100111001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100100111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100101000010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000100101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000100101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1000100101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000100110001000" => 
 	 	 	 	 color <= "110001";
 	 	 	when "1000100110001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100110001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100110001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100110001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100110001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100110001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000100110001111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "1000100110010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000100110010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000100110010010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1000100110010011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000100110010100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000101000111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101000111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101001000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101001000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101001000010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000101001000011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000101001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000101001101011" => 
 	 	 	 	 color <= "101111";
 	 	 	when "1000101001101100" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1000101001101101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1000101001101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1000101001101111" => 
 	 	 	 	 color <= "011010";
 	 	 	when "1000101001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000101010000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000101010001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101010001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101010001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101010001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101010001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101010001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101010001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101010001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101010010000" => 
 	 	 	 	 color <= "111010";
 	 	 	when "1000101010010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000101010010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000101010010011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000101010010100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000101010010101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1000101100111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101100111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101100111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101100111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101100111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101101000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101101000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101101000010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000101101000011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000101101101010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1000101101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000101101101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000101101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000101101101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000101101101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000101101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000101110000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101110001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101110001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101110001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101110001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101110001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101110001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101110001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101110001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101110010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000101110010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000101110010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000101110010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000101110010100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000101110010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000110000111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110000111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110000111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110000111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110001000000" => 
 	 	 	 	 color <= "100101";
 	 	 	when "1000110001000001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000110001000010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000110001000011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000110001101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000110001101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000110001101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000110001101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000110001101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000110001110000" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1000110010000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1000110010000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110010001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110010001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110010001010" => 
 	 	 	 	 color <= "110001";
 	 	 	when "1000110010001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1000110010001100" => 
 	 	 	 	 color <= "110001";
 	 	 	when "1000110010001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110010001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110010001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110010010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110010010001" => 
 	 	 	 	 color <= "111010";
 	 	 	when "1000110010010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000110010010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000110010010100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000110010010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000110010010110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1000110100111101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000110100111110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000110100111111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000110101000000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000110101000001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000110101000010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000110101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000110101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000110101101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000110101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000110101101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000110101101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000110101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000110110000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110110000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110110001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110110001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110110001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1000110110001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110110001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110110001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110110010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110110010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000110110010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000110110010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000110110010100" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1000110110010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000110110010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000111000111111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000111001000000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000111001101010" => 
 	 	 	 	 color <= "010001";
 	 	 	when "1000111001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000111001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000111001101101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1000111001101110" => 
 	 	 	 	 color <= "010001";
 	 	 	when "1000111001101111" => 
 	 	 	 	 color <= "010001";
 	 	 	when "1000111001110000" => 
 	 	 	 	 color <= "010001";
 	 	 	when "1000111010000101" => 
 	 	 	 	 color <= "100001";
 	 	 	when "1000111010000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111010000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111010001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111010001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111010001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111010001011" => 
 	 	 	 	 color <= "110001";
 	 	 	when "1000111010001100" => 
 	 	 	 	 color <= "110001";
 	 	 	when "1000111010001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111010001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111010001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111010010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111010010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111010010010" => 
 	 	 	 	 color <= "111010";
 	 	 	when "1000111010010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000111010010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000111010010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000111010010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000111101101011" => 
 	 	 	 	 color <= "010001";
 	 	 	when "1000111101101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000111101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1000111110000100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1000111110000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111110000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111110000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111110001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111110001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111110001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111110001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111110001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111110001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111110001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111110001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111110010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111110010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1000111110010010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "1000111110010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000111110010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1000111110010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000111110010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1000111110010111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1001000001101100" => 
 	 	 	 	 color <= "010001";
 	 	 	when "1001000001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001000001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001000010000100" => 
 	 	 	 	 color <= "110001";
 	 	 	when "1001000010000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000010000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000010000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000010001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000010001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000010001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000010001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000010001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000010001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000010001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000010001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000010010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000010010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000010010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000010010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001000010010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001000010010101" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1001000010010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001000010010111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1001000101101101" => 
 	 	 	 	 color <= "010001";
 	 	 	when "1001000101101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001000101101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001000110000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1001000110000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000110000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000110000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000110000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000110001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000110001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000110001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000110001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000110001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1001000110001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000110001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000110001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000110010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000110010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000110010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001000110010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001000110010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001000110010101" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1001000110010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001000110010111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1001001001101010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1001001001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1001001001101100" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1001001001101101" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1001001001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001001001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001001001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001001010000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001010000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001010000101" => 
 	 	 	 	 color <= "100001";
 	 	 	when "1001001010000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1001001010001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001010001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001010001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001010001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001010001101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1001001010001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001010001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001010010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001010010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001010010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001010010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001001010010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001001010010101" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1001001010010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001001010010111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1001001101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001001101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001001101101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001001101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001001101101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001001101101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001001101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001001110000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1001001110000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001110000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001110000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001110000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1001001110000111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1001001110001000" => 
 	 	 	 	 color <= "110001";
 	 	 	when "1001001110001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001110001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001110001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001110001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1001001110001101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1001001110001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001110001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001110010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001110010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001110010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001001110010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001001110010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001001110010101" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1001001110010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001001110010111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001010010000001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1001010010000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010010010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001010010010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001010010010101" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1001010010010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001010010010111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1001010110000001" => 
 	 	 	 	 color <= "110001";
 	 	 	when "1001010110000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001010110010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001010110010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001010110010101" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1001010110010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001010110010111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1001011010000000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1001011010000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011010000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011010000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011010000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011010000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011010000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011010000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011010001000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1001011010001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1001011010001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011010001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011010001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011010001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011010001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011010001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011010010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011010010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011010010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011010010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001011010010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001011010010101" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1001011010010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001011010010111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1001011110000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110001000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1001011110001001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1001011110001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001011110010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001011110010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001011110010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001011110010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001011110010111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1001100001101010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1001100001101011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1001100001111111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1001100010000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100010000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100010000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100010000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100010000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100010000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100010000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100010000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100010001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1001100010001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1001100010001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100010001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100010001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100010001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100010001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100010001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100010010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100010010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100010010010" => 
 	 	 	 	 color <= "111010";
 	 	 	when "1001100010010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001100010010100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001100010010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001100010010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001100101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001100101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1001100101111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100110000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100110000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100110000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100110000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100110000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100110000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100110000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100110000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100110001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100110001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100110001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100110001011" => 
 	 	 	 	 color <= "110001";
 	 	 	when "1001100110001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1001100110001101" => 
 	 	 	 	 color <= "110001";
 	 	 	when "1001100110001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100110001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100110010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100110010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001100110010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001100110010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001100110010100" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1001100110010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001100110010110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001101001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001101001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1001101001111110" => 
 	 	 	 	 color <= "100001";
 	 	 	when "1001101001111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101010000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101010000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101010000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101010000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101010000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101010000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1001101010000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1001101010000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101010001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101010001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101010001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101010001011" => 
 	 	 	 	 color <= "100001";
 	 	 	when "1001101010001110" => 
 	 	 	 	 color <= "110001";
 	 	 	when "1001101010001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101010010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101010010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101010010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001101010010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001101010010100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001101010010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001101010010110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1001101101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001101101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001101101101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001101101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001101101101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001101101101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001101101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001101101111101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1001101101111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101101111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101110000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101110000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101110000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101110000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101110000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101110000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1001101110000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101110001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101110001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101110001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101110001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101110001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101110001101" => 
 	 	 	 	 color <= "110001";
 	 	 	when "1001101110001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101110001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101110010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001101110010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001101110010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001101110010011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001101110010100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001101110010101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001110001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001110001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001110001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001110001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001110001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001110001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001110001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001110001111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110001111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110001111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110010000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110010000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110010000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110010000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110010000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110010000101" => 
 	 	 	 	 color <= "110001";
 	 	 	when "1001110010000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1001110010000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110010001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110010001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110010001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110010001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110010001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110010001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110010001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110010001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110010010000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "1001110010010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001110010010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001110010010011" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1001110010010100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001110010010101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1001110100101010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1001110100101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001110100101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001110100101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001110100101110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1001110101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001110101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1001110101111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1001110101111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110101111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110101111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110001111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001110110010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001110110010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001110110010010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001110110010011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001110110010100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001111000101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111000101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111000101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111000101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111000101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111000101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111000101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111000101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111000110000" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1001111001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1001111001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1001111001111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111001111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111001111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111001111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111010000000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1001111010000001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1001111010000010" => 
 	 	 	 	 color <= "110001";
 	 	 	when "1001111010000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111010000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111010000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111010000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111010000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111010001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111010001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111010001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111010001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111010001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111010001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111010001110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111010001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001111010010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001111010010001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001111010010010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001111010010011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001111010010100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1001111100100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111100101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111100101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111100101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111100101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111100101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111100101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111100101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111100101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111100110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111100110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111101101010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1001111101101011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1001111101111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1001111101111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111101111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111101111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111101111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111110000000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1001111110000001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1001111110000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1001111110000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111110000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111110000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111110000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111110000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111110001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111110001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111110001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111110001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111110001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111110001101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1001111110001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001111110001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001111110010000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1001111110010001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1001111110010010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1001111110010011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010000000100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000000100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000000101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000000101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000000101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000000101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000000101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000000101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000000101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000000101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000000110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000000110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000000110010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010000001101010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1010000001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010000001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010000001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010000001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010000001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010000001110000" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1010000001111010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1010000001111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000001111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000001111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000001111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000001111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000010000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000010000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000010000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000010000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000010000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000010000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1010000010000110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1010000010000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000010001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000010001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000010001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000010001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000010001100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000010001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010000010001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010000010001111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010000010010000" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010000010010001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010000010010010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010000100100101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010000100100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000100100111" => 
 	 	 	 	 color <= "000110";
 	 	 	when "1010000100101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000100101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000100101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000100101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000100101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000100101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000100101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000100101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000100110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000100110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000100110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010000101101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010000101101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010000101101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010000101101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010000101101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010000101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010000101111010" => 
 	 	 	 	 color <= "110001";
 	 	 	when "1010000101111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000101111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000101111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000101111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000101111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000110000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000110000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000110000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000110000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000110000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000110000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "1010000110000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000110001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000110001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000110001010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000110001011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010000110001100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010000110001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010000110001110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010000110001111" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010000110010000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010000110010001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010000110010010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1010001000100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001000100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001000100111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010001000101000" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010001000101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001000101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001000101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001000101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001000101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001000101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001000101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001000110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001000110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001000110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001000110011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010001001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010001001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1010001001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010001001111001" => 
 	 	 	 	 color <= "100101";
 	 	 	when "1010001001111010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001001111011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001001111100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001001111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001001111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001001111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001010000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001010000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001010000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001010000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001010000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001010000101" => 
 	 	 	 	 color <= "110001";
 	 	 	when "1010001010000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "1010001010000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001010001000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001010001001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001010001010" => 
 	 	 	 	 color <= "111010";
 	 	 	when "1010001010001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010001010001100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010001010001101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010001010001110" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010001010001111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010001010010000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010001010010001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1010001100011101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1010001100011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010001100011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010001100100000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010001100100001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1010001100100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001100100110" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010001100100111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010001100101000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010001100101001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010001100101010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010001100101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001100101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001100101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001100101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001100101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001100110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001100110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001100110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001100110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010001101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1010001101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010001101111001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010001101111010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010001101111011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010001101111100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "1010001101111101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001101111110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001101111111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001110000000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001110000001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001110000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001110000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001110000100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001110000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001110000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001110000111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "1010001110001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010001110001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010001110001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010001110001011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010001110001100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010001110001101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010001110001110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010001110001111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010001110010000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1010010000011101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1010010000011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010000011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010000100000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010000100001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010000100010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010000100011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010000100100" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1010010000100101" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010010000100110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010010000100111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010010000101000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010010000101001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010010000101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010000101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010000101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010000101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010000101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010000101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010000110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010000110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010000110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010000110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010001101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010010001101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1010010001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010010001111000" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1010010001111001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010001111010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010001111011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010001111100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010001111101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010001111110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010001111111" => 
 	 	 	 	 color <= "111010";
 	 	 	when "1010010010000000" => 
 	 	 	 	 color <= "111010";
 	 	 	when "1010010010000001" => 
 	 	 	 	 color <= "111010";
 	 	 	when "1010010010000010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "1010010010000011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "1010010010000100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "1010010010000101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010010000110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010010000111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010010001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010010001001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010010001010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010010001011" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010010010001100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010010001101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010010001110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010010001111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1010010100011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010100011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010100100000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010100100001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010100100010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010100100011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010100100100" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1010010100100101" => 
 	 	 	 	 color <= "000110";
 	 	 	when "1010010100100110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010010100100111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010010100101000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010010100101001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010010100101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010100101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010100101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010100101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010100101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010100101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010100110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010100110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010100110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010100110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010101101010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010010101101011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "1010010101101111" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010010101110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010010101111000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010101111001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010101111010" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010010101111011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010101111100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010101111101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010101111110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010101111111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010110000000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010110000001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010110000010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010110000011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010110000100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010110000101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010110000110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010110000111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010110001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010010110001001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010010110001010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010110001011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010110001100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010010110001101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011000011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011000011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011000100000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011000100001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011000100010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011000100011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011000100100" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1010011000100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011000100110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010011000100111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010011000101000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010011000101001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010011000101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011000101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011000101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011000101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011000101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011000101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011000110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011000110001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010011000110010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010011000110011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010011001101010" => 
 	 	 	 	 color <= "111011";
 	 	 	when "1010011001101011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010011001101100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010011001101101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010011001101110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010011001101111" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010011001110000" => 
 	 	 	 	 color <= "111111";
 	 	 	when "1010011001111000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011001111001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011001111010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011001111011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011001111100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011001111101" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010011001111110" => 
 	 	 	 	 color <= "101110";
 	 	 	when "1010011001111111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010011010000000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010011010000001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010011010000010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010011010000011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010011010000100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "1010011010000101" => 
 	 	 	 	 color <= "101110";
 	 	 	when "1010011010000110" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010011010000111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011010001000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011010001001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011010001010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011010001011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011010001100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1010011100011110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1010011100011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011100100000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011100100001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011100100010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011100100011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011100100100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011100100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011100100110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010011100100111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010011100101000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010011100101001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010011100101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011100101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011100101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011100101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011100101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011100101111" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010011100110000" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010011100110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011100110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011100110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011100110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011100110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011100110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011100110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011101101011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1010011101101100" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1010011101101101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1010011101101110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1010011101101111" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1010011101111001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1010011101111010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011101111011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011101111100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011101111101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011101111110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011101111111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011110000000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011110000001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011110000010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011110000011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011110000100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011110000101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011110000110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011110000111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011110001000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011110001001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010011110001010" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1010100000011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100000100000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100000100001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100000100010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100000100011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100000100100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100000100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100000100110" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010100000100111" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010100000101000" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010100000101001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010100000101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100000101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100000101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100000101101" => 
 	 	 	 	 color <= "000110";
 	 	 	when "1010100000101110" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010100000101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100000110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100000110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100000110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100000110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100000110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100000110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100000110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100000110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100000111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100000111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100001111100" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1010100001111101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1010100001111110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100001111111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100010000000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100010000001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100010000010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100010000011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100010000100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100010000101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100010000110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1010100010000111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "1010100100011111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1010100100100000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100100100001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100100100010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100100100011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100100100100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010100100100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100101101" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010100100101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000100000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1010101000100001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010101000100010" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010101000100011" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010101000100100" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010101000100101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010101000100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000101100" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010101000101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100100000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010101100100001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010101100100010" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010101100100011" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010101100100100" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010101100100101" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010101100100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100101011" => 
 	 	 	 	 color <= "000110";
 	 	 	when "1010101100101100" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010101100101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100111100" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010110000011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010110000100000" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010110000100001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010110000100010" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010110000100011" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010110000100100" => 
 	 	 	 	 color <= "011010";
 	 	 	when "1010110000100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000100110" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010110000100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000101011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010110000101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000101111" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010110000110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100011110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "1010110100011111" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010110100100000" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010110100100001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010110100100010" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010110100100011" => 
 	 	 	 	 color <= "011010";
 	 	 	when "1010110100100100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100100110" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010110100100111" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010110100101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100101011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010110100101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100101111" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010110100110000" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010110100110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100111101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010111000011110" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010111000011111" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010111000100000" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010111000100001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010111000100010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1010111000100011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111000100100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111000100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111000100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111000100111" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010111000101000" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010111000101001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010111000101010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010111000101011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010111000101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111000101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111000101110" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010111000101111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010111000110000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010111000110001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010111000110010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010111000110011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010111000110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111000110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111000110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111000110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111000111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111000111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111000111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111000111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111000111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111000111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100011101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1010111100011110" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010111100011111" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010111100100000" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010111100100001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "1010111100100010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100100011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100100100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100101001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010111100101010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010111100101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100101110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010111100101111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010111100110000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010111100110001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1010111100110010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010111100110011" => 
 	 	 	 	 color <= "000110";
 	 	 	when "1010111100110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000011101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "1011000000011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1011000000011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1011000000100000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1011000000100001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "1011000000100010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000100011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000100100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000101010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011000000101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000101101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011000000101110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011000000101111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011000000110000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011000000110001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011000000110010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011000000110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000000111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100100001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011000100100010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100100011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100100100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100101010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011000100101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100101101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011000100101110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011000100101111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011000100110000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011000100110001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011000100110010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011000100110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000100001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011001000100010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000100011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000100100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000101010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011001000101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000101110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011001000101111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011001000110000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011001000110001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011001000110010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011001000110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100100001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011001100100010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100100011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011001100100100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011001100100101" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011001100100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100101010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011001100101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100101110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011001100101111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011001100110000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011001100110001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011001100110010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011001100110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000100010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000100011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011010000100100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011010000100101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011010000100110" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011010000100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000101010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011010000101011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011010000101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000101110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011010000101111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011010000110000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011010000110001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011010000110010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011010000110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000111101" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011010100100010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100100011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011010100100100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011010100100101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011010100100110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011010100100111" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011010100101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100101011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011010100101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100101110" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011010100101111" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011010100110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000100011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000100100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011011000100101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011011000100110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011011000100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000101011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011011000101100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011011000101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100100011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011011100100100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100100110" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011011100100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100101011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011011100101101" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011011100101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100000111011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011100100101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100100110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100100110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100100110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100100110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100100110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100100110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100100110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100100110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100100111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100100111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101000110000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011101000110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101000110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101000110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101000110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101000110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101000110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101000110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101000111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101100110011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011101100110100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011101100110101" => 
 	 	 	 	 color <= "000001"; 
 	 	 end case; 
     	 end if;  
     end process; 
 address <= row & col; 
 end;
