library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ROM is
  port(
	  row : in std_logic_vector(4 downto 0);
	  col : in std_logic_vector(4 downto 0);
	  fruit_color : in std_logic_vector(5 downto 0);
	  clk : in std_logic;
	  color : out std_logic_vector(5 downto 0)
  );
end ROM;

architecture synth of ROM is 
signal address : std_logic_vector(9 downto 0);
begin
	process(clk) is
	begin
		if rising_edge(clk) then
			case address is 

 	 	 	when 0000001100=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000001101=> 
 	 	 	 	 <= GFGFGD
 	 	 	when 0000001110=> 
 	 	 	 	 <= GFG4F3
 	 	 	when 0000001111=> 
 	 	 	 	 <= GEFFE3
 	 	 	when 0000010000=> 
 	 	 	 	 <= GEFEE1
 	 	 	when 0000010001=> 
 	 	 	 	 <= GFG2EG
 	 	 	when 0000010010=> 
 	 	 	 	 <= GFGEGB
 	 	 	when 0000010011=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000101001=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000101010=> 
 	 	 	 	 <= GEF7D1
 	 	 	when 0000101011=> 
 	 	 	 	 <= GCD66C
 	 	 	when 0000101100=> 
 	 	 	 	 <= G9BD28
 	 	 	when 0000101101=> 
 	 	 	 	 <= G99E01
 	 	 	when 0000101110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0000101111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0000110000=> 
 	 	 	 	 <= G89D00
 	 	 	when 0000110001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0000110010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0000110011=> 
 	 	 	 	 <= G9B81G
 	 	 	when 0000110100=> 
 	 	 	 	 <= GCD15G
 	 	 	when 0000110101=> 
 	 	 	 	 <= GEF1C2
 	 	 	when 0000110110=> 
 	 	 	 	 <= GFGEGC
 	 	 	when 0001000111=> 
 	 	 	 	 <= GFGFGE
 	 	 	when 0001001000=> 
 	 	 	 	 <= GDE89D
 	 	 	when 0001001001=> 
 	 	 	 	 <= G9B91G
 	 	 	when 0001001010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0001001011=> 
 	 	 	 	 <= G99E01
 	 	 	when 0001001100=> 
 	 	 	 	 <= GBBE26
 	 	 	when 0001001101=> 
 	 	 	 	 <= GCCG50
 	 	 	when 0001001110=> 
 	 	 	 	 <= GDDC6C
 	 	 	when 0001001111=> 
 	 	 	 	 <= GDE179
 	 	 	when 0001010000=> 
 	 	 	 	 <= GDE178
 	 	 	when 0001010001=> 
 	 	 	 	 <= GDDD6D
 	 	 	when 0001010010=> 
 	 	 	 	 <= GCD051
 	 	 	when 0001010011=> 
 	 	 	 	 <= GBBF28
 	 	 	when 0001010100=> 
 	 	 	 	 <= G99E01
 	 	 	when 0001010101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0001010110=> 
 	 	 	 	 <= G9B312
 	 	 	when 0001010111=> 
 	 	 	 	 <= GDDG84
 	 	 	when 0001011000=> 
 	 	 	 	 <= GFGCG6
 	 	 	when 0001100101=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0001100110=> 
 	 	 	 	 <= GEFEE0
 	 	 	when 0001100111=> 
 	 	 	 	 <= G9BD29
 	 	 	when 0001101000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0001101001=> 
 	 	 	 	 <= G9B719
 	 	 	when 0001101010=> 
 	 	 	 	 <= GDDE70
 	 	 	when 0001101011=> 
 	 	 	 	 <= GFFCC5
 	 	 	when 0001101100=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0001101101=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0001101110=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 0001101111=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0001110000=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0001110001=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0001110010=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0001110011=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0001110100=> 
 	 	 	 	 <= GFFDC7
 	 	 	when 0001110101=> 
 	 	 	 	 <= GDDG74
 	 	 	when 0001110110=> 
 	 	 	 	 <= G9B91E
 	 	 	when 0001110111=> 
 	 	 	 	 <= G99D00
 	 	 	when 0001111000=> 
 	 	 	 	 <= G9B516
 	 	 	when 0001111001=> 
 	 	 	 	 <= GEF2C4
 	 	 	when 0010000100=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0010000101=> 
 	 	 	 	 <= GDE89B
 	 	 	when 0010000110=> 
 	 	 	 	 <= G99F03
 	 	 	when 0010000111=> 
 	 	 	 	 <= G9B008
 	 	 	when 0010001000=> 
 	 	 	 	 <= GDDG73
 	 	 	when 0010001001=> 
 	 	 	 	 <= GFG0CG
 	 	 	when 0010001010=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 0010001011=> 
 	 	 	 	 <= GFF9BG
 	 	 	when 0010001100=> 
 	 	 	 	 <= GDDE70
 	 	 	when 0010001101=> 
 	 	 	 	 <= GBC83G
 	 	 	when 0010001110=> 
 	 	 	 	 <= GBBB1G
 	 	 	when 0010001111=> 
 	 	 	 	 <= G9B410
 	 	 	when 0010010000=> 
 	 	 	 	 <= GBBD22
 	 	 	when 0010010001=> 
 	 	 	 	 <= GCC941
 	 	 	when 0010010010=> 
 	 	 	 	 <= GFFEC9
 	 	 	when 0010010011=> 
 	 	 	 	 <= GFF7BD
 	 	 	when 0010010100=> 
 	 	 	 	 <= GFF8BF
 	 	 	when 0010010101=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0010010110=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0010010111=> 
 	 	 	 	 <= GDE27B
 	 	 	when 0010011000=> 
 	 	 	 	 <= G9B20D
 	 	 	when 0010011001=> 
 	 	 	 	 <= G99D00
 	 	 	when 0010011010=> 
 	 	 	 	 <= GCD871
 	 	 	when 0010011011=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0010100011=> 
 	 	 	 	 <= GFGFGG
 	 	 	when 0010100100=> 
 	 	 	 	 <= GDDF82
 	 	 	when 0010100101=> 
 	 	 	 	 <= G99D00
 	 	 	when 0010100110=> 
 	 	 	 	 <= GBBD24
 	 	 	when 0010100111=> 
 	 	 	 	 <= GFF7BC
 	 	 	when 0010101000=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0010101001=> 
 	 	 	 	 <= GFFFCB
 	 	 	when 0010101010=> 
 	 	 	 	 <= GBC83G
 	 	 	when 0010101011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0010101100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0010101101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0010101110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0010101111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0010110000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0010110001=> 
 	 	 	 	 <= G99D00
 	 	 	when 0010110010=> 
 	 	 	 	 <= GFFCC4
 	 	 	when 0010110011=> 
 	 	 	 	 <= G99G06
 	 	 	when 0010110100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0010110101=> 
 	 	 	 	 <= GBC537
 	 	 	when 0010110110=> 
 	 	 	 	 <= GEF29G
 	 	 	when 0010110111=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0010111000=> 
 	 	 	 	 <= GFFBC1
 	 	 	when 0010111001=> 
 	 	 	 	 <= GBBG2C
 	 	 	when 0010111010=> 
 	 	 	 	 <= G89D00
 	 	 	when 0010111011=> 
 	 	 	 	 <= GCCF58
 	 	 	when 0010111100=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0011000011=> 
 	 	 	 	 <= GDE798
 	 	 	when 0011000100=> 
 	 	 	 	 <= G99D00
 	 	 	when 0011000101=> 
 	 	 	 	 <= GBC130
 	 	 	when 0011000110=> 
 	 	 	 	 <= GFFFCC
 	 	 	when 0011000111=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0011001000=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0011001001=> 
 	 	 	 	 <= GEEB8E
 	 	 	when 0011001010=> 
 	 	 	 	 <= G99D00
 	 	 	when 0011001011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011001100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011001101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011001110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011001111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011010000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011010001=> 
 	 	 	 	 <= G9B719
 	 	 	when 0011010010=> 
 	 	 	 	 <= GEF09B
 	 	 	when 0011010011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011010100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011010101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011010110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011010111=> 
 	 	 	 	 <= GCD45B
 	 	 	when 0011011000=> 
 	 	 	 	 <= GFG0CG
 	 	 	when 0011011001=> 
 	 	 	 	 <= GFFGCE
 	 	 	when 0011011010=> 
 	 	 	 	 <= GBC537
 	 	 	when 0011011011=> 
 	 	 	 	 <= G99D00
 	 	 	when 0011011100=> 
 	 	 	 	 <= GCD76E
 	 	 	when 0011011101=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0011100010=> 
 	 	 	 	 <= GEFDDG
 	 	 	when 0011100011=> 
 	 	 	 	 <= G99F03
 	 	 	when 0011100100=> 
 	 	 	 	 <= GBBC21
 	 	 	when 0011100101=> 
 	 	 	 	 <= GFFFCB
 	 	 	when 0011100110=> 
 	 	 	 	 <= GFG0CG
 	 	 	when 0011100111=> 
 	 	 	 	 <= GCD358
 	 	 	when 0011101000=> 
 	 	 	 	 <= GBC334
 	 	 	when 0011101001=> 
 	 	 	 	 <= GFF3B2
 	 	 	when 0011101010=> 
 	 	 	 	 <= GBC437
 	 	 	when 0011101011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011101100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011101101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011101110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011101111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011110000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011110001=> 
 	 	 	 	 <= GCCD48
 	 	 	when 0011110010=> 
 	 	 	 	 <= GDDC6D
 	 	 	when 0011110011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011110100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011110101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011110110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011110111=> 
 	 	 	 	 <= G99D00
 	 	 	when 0011111000=> 
 	 	 	 	 <= GBC538
 	 	 	when 0011111001=> 
 	 	 	 	 <= GFG0CG
 	 	 	when 0011111010=> 
 	 	 	 	 <= GFFFCD
 	 	 	when 0011111011=> 
 	 	 	 	 <= GBBE26
 	 	 	when 0011111100=> 
 	 	 	 	 <= G89D00
 	 	 	when 0011111101=> 
 	 	 	 	 <= GEEFB9
 	 	 	when 0100000001=> 
 	 	 	 	 <= GFGFGE
 	 	 	when 0100000010=> 
 	 	 	 	 <= GBBE2C
 	 	 	when 0100000011=> 
 	 	 	 	 <= G99G05
 	 	 	when 0100000100=> 
 	 	 	 	 <= GFF6B8
 	 	 	when 0100000101=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0100000110=> 
 	 	 	 	 <= GCCB43
 	 	 	when 0100000111=> 
 	 	 	 	 <= G89D00
 	 	 	when 0100001000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100001001=> 
 	 	 	 	 <= G9B616
 	 	 	when 0100001010=> 
 	 	 	 	 <= GFF8BD
 	 	 	when 0100001011=> 
 	 	 	 	 <= G9B616
 	 	 	when 0100001100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100001101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100001110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100001111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100010000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100010001=> 
 	 	 	 	 <= GDE077
 	 	 	when 0100010010=> 
 	 	 	 	 <= GBC73E
 	 	 	when 0100010011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100010100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100010101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100010110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100010111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100011000=> 
 	 	 	 	 <= G99D00
 	 	 	when 0100011001=> 
 	 	 	 	 <= GFF6B8
 	 	 	when 0100011010=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0100011011=> 
 	 	 	 	 <= GFF8BE
 	 	 	when 0100011100=> 
 	 	 	 	 <= G9B008
 	 	 	when 0100011101=> 
 	 	 	 	 <= G9B30G
 	 	 	when 0100011110=> 
 	 	 	 	 <= GFG9G1
 	 	 	when 0100100001=> 
 	 	 	 	 <= GDEDB4
 	 	 	when 0100100010=> 
 	 	 	 	 <= G99D00
 	 	 	when 0100100011=> 
 	 	 	 	 <= GDD863
 	 	 	when 0100100100=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0100100101=> 
 	 	 	 	 <= GDE076
 	 	 	when 0100100110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100100111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100101000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100101001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100101010=> 
 	 	 	 	 <= GBC538
 	 	 	when 0100101011=> 
 	 	 	 	 <= GEF19F
 	 	 	when 0100101100=> 
 	 	 	 	 <= G99F04
 	 	 	when 0100101101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100101110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100101111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100110000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100110001=> 
 	 	 	 	 <= GFF5B5
 	 	 	when 0100110010=> 
 	 	 	 	 <= G9B30G
 	 	 	when 0100110011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100110100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100110101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100110110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100110111=> 
 	 	 	 	 <= G9B20D
 	 	 	when 0100111000=> 
 	 	 	 	 <= GEE47G
 	 	 	when 0100111001=> 
 	 	 	 	 <= GFF6B9
 	 	 	when 0100111010=> 
 	 	 	 	 <= GFFDC7
 	 	 	when 0100111011=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0100111100=> 
 	 	 	 	 <= GDDD6E
 	 	 	when 0100111101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100111110=> 
 	 	 	 	 <= GCDB76
 	 	 	when 0101000000=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0101000001=> 
 	 	 	 	 <= GBBF2D
 	 	 	when 0101000010=> 
 	 	 	 	 <= G9B009
 	 	 	when 0101000011=> 
 	 	 	 	 <= GFFFCB
 	 	 	when 0101000100=> 
 	 	 	 	 <= GFFEC9
 	 	 	when 0101000101=> 
 	 	 	 	 <= G9B10B
 	 	 	when 0101000110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101000111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101001000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101001001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101001010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101001011=> 
 	 	 	 	 <= GDD965
 	 	 	when 0101001100=> 
 	 	 	 	 <= GDE077
 	 	 	when 0101001101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101001110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101001111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101010000=> 
 	 	 	 	 <= G9B109
 	 	 	when 0101010001=> 
 	 	 	 	 <= GFF8BE
 	 	 	when 0101010010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101010011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101010100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101010101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101010110=> 
 	 	 	 	 <= GCC840
 	 	 	when 0101010111=> 
 	 	 	 	 <= GFF7BC
 	 	 	when 0101011000=> 
 	 	 	 	 <= GCCE4C
 	 	 	when 0101011001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101011010=> 
 	 	 	 	 <= G9B007
 	 	 	when 0101011011=> 
 	 	 	 	 <= GFFBC2
 	 	 	when 0101011100=> 
 	 	 	 	 <= GFFGCE
 	 	 	when 0101011101=> 
 	 	 	 	 <= G9B30G
 	 	 	when 0101011110=> 
 	 	 	 	 <= G9B10C
 	 	 	when 0101100000=> 
 	 	 	 	 <= GFG1EC
 	 	 	when 0101100001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101100010=> 
 	 	 	 	 <= GCCG4G
 	 	 	when 0101100011=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0101100100=> 
 	 	 	 	 <= GEF2B0
 	 	 	when 0101100101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101100110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101100111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101101000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101101001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101101010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101101011=> 
 	 	 	 	 <= G99E01
 	 	 	when 0101101100=> 
 	 	 	 	 <= GEEC90
 	 	 	when 0101101101=> 
 	 	 	 	 <= GCCD48
 	 	 	when 0101101110=> 
 	 	 	 	 <= G89D00
 	 	 	when 0101101111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101110000=> 
 	 	 	 	 <= GBC435
 	 	 	when 0101110001=> 
 	 	 	 	 <= GEE37F
 	 	 	when 0101110010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101110011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101110100=> 
 	 	 	 	 <= G9B310
 	 	 	when 0101110101=> 
 	 	 	 	 <= GEE786
 	 	 	when 0101110110=> 
 	 	 	 	 <= GEE98B
 	 	 	when 0101110111=> 
 	 	 	 	 <= G9B412
 	 	 	when 0101111000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101111001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101111010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101111011=> 
 	 	 	 	 <= GCD55D
 	 	 	when 0101111100=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0101111101=> 
 	 	 	 	 <= GCD45B
 	 	 	when 0101111110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110000000=> 
 	 	 	 	 <= GDE490
 	 	 	when 0110000001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110000010=> 
 	 	 	 	 <= GEEB8E
 	 	 	when 0110000011=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0110000100=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0110000101=> 
 	 	 	 	 <= GCD55F
 	 	 	when 0110000110=> 
 	 	 	 	 <= G9B717
 	 	 	when 0110000111=> 
 	 	 	 	 <= G99D00
 	 	 	when 0110001000=> 
 	 	 	 	 <= G89D00
 	 	 	when 0110001001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110001010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110001011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110001100=> 
 	 	 	 	 <= G9B20E
 	 	 	when 0110001101=> 
 	 	 	 	 <= GFF7BB
 	 	 	when 0110001110=> 
 	 	 	 	 <= GBBC21
 	 	 	when 0110001111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110010000=> 
 	 	 	 	 <= GDD864
 	 	 	when 0110010001=> 
 	 	 	 	 <= GCCG4G
 	 	 	when 0110010010=> 
 	 	 	 	 <= G89D00
 	 	 	when 0110010011=> 
 	 	 	 	 <= GCCC47
 	 	 	when 0110010100=> 
 	 	 	 	 <= GFF7BC
 	 	 	when 0110010101=> 
 	 	 	 	 <= GCCB44
 	 	 	when 0110010110=> 
 	 	 	 	 <= G99D00
 	 	 	when 0110010111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110011000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110011001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110011010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110011011=> 
 	 	 	 	 <= G9B513
 	 	 	when 0110011100=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0110011101=> 
 	 	 	 	 <= GEEG99
 	 	 	when 0110011110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110100000=> 
 	 	 	 	 <= GCCG5B
 	 	 	when 0110100001=> 
 	 	 	 	 <= G99D00
 	 	 	when 0110100010=> 
 	 	 	 	 <= GFFEC9
 	 	 	when 0110100011=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0110100100=> 
 	 	 	 	 <= GEEF96
 	 	 	when 0110100101=> 
 	 	 	 	 <= GDE37E
 	 	 	when 0110100110=> 
 	 	 	 	 <= GEED93
 	 	 	when 0110100111=> 
 	 	 	 	 <= GFF9C0
 	 	 	when 0110101000=> 
 	 	 	 	 <= GEEC90
 	 	 	when 0110101001=> 
 	 	 	 	 <= GDD967
 	 	 	when 0110101010=> 
 	 	 	 	 <= GBC73F
 	 	 	when 0110101011=> 
 	 	 	 	 <= G9B514
 	 	 	when 0110101100=> 
 	 	 	 	 <= G99D00
 	 	 	when 0110101101=> 
 	 	 	 	 <= GBBG2C
 	 	 	when 0110101110=> 
 	 	 	 	 <= GFF7BC
 	 	 	when 0110101111=> 
 	 	 	 	 <= GBC334
 	 	 	when 0110110000=> 
 	 	 	 	 <= GFF7BB
 	 	 	when 0110110001=> 
 	 	 	 	 <= GBC83F
 	 	 	when 0110110010=> 
 	 	 	 	 <= GEEB8E
 	 	 	when 0110110011=> 
 	 	 	 	 <= GEE684
 	 	 	when 0110110100=> 
 	 	 	 	 <= G9B30F
 	 	 	when 0110110101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110110110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110110111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110111000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110111001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110111010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110111011=> 
 	 	 	 	 <= G99D00
 	 	 	when 0110111100=> 
 	 	 	 	 <= GFF8BD
 	 	 	when 0110111101=> 
 	 	 	 	 <= GFG0CF
 	 	 	when 0110111110=> 
 	 	 	 	 <= G99E01
 	 	 	when 0111000000=> 
 	 	 	 	 <= GBC238
 	 	 	when 0111000001=> 
 	 	 	 	 <= G9B009
 	 	 	when 0111000010=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0111000011=> 
 	 	 	 	 <= GFF5B7
 	 	 	when 0111000100=> 
 	 	 	 	 <= G99E01
 	 	 	when 0111000101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111000110=> 
 	 	 	 	 <= G99D00
 	 	 	when 0111000111=> 
 	 	 	 	 <= G99D00
 	 	 	when 0111001000=> 
 	 	 	 	 <= G9B718
 	 	 	when 0111001001=> 
 	 	 	 	 <= GCC941
 	 	 	when 0111001010=> 
 	 	 	 	 <= GDDC6B
 	 	 	when 0111001011=> 
 	 	 	 	 <= GEEE94
 	 	 	when 0111001100=> 
 	 	 	 	 <= GFF9BG
 	 	 	when 0111001101=> 
 	 	 	 	 <= GFF2B0
 	 	 	when 0111001110=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0111001111=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0111010000=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0111010001=> 
 	 	 	 	 <= GFFEC8
 	 	 	when 0111010010=> 
 	 	 	 	 <= GBC73E
 	 	 	when 0111010011=> 
 	 	 	 	 <= G89D00
 	 	 	when 0111010100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111010101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111010110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111010111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111011000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111011001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111011010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111011011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111011100=> 
 	 	 	 	 <= GEEB8E
 	 	 	when 0111011101=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0111011110=> 
 	 	 	 	 <= G9B514
 	 	 	when 0111100000=> 
 	 	 	 	 <= GBBE2B
 	 	 	when 0111100001=> 
 	 	 	 	 <= G9B513
 	 	 	when 0111100010=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0111100011=> 
 	 	 	 	 <= GEE98D
 	 	 	when 0111100100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111100101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111100110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111100111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111101000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111101001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111101010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111101011=> 
 	 	 	 	 <= G99D00
 	 	 	when 0111101100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111101101=> 
 	 	 	 	 <= GCCC47
 	 	 	when 0111101110=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0111101111=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0111110000=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0111110001=> 
 	 	 	 	 <= GFFGCE
 	 	 	when 0111110010=> 
 	 	 	 	 <= GEEB8E
 	 	 	when 0111110011=> 
 	 	 	 	 <= GDD863
 	 	 	when 0111110100=> 
 	 	 	 	 <= GBC63B
 	 	 	when 0111110101=> 
 	 	 	 	 <= G9B411
 	 	 	when 0111110110=> 
 	 	 	 	 <= G99D00
 	 	 	when 0111110111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111111000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111111001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111111010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111111011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111111100=> 
 	 	 	 	 <= GEE887
 	 	 	when 0111111101=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0111111110=> 
 	 	 	 	 <= G9B91E
 	 	 	when 1000000000=> 
 	 	 	 	 <= GBBG2G
 	 	 	when 1000000001=> 
 	 	 	 	 <= G9B30F
 	 	 	when 1000000010=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1000000011=> 
 	 	 	 	 <= GEEC90
 	 	 	when 1000000100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000000101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000000110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000000111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000001000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000001001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000001010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000001011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000001100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000001101=> 
 	 	 	 	 <= GDE27C
 	 	 	when 1000001110=> 
 	 	 	 	 <= GFFEC8
 	 	 	when 1000001111=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1000010000=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1000010001=> 
 	 	 	 	 <= GDD863
 	 	 	when 1000010010=> 
 	 	 	 	 <= GBBB20
 	 	 	when 1000010011=> 
 	 	 	 	 <= GCCB45
 	 	 	when 1000010100=> 
 	 	 	 	 <= GDDD6F
 	 	 	when 1000010101=> 
 	 	 	 	 <= GEEF97
 	 	 	when 1000010110=> 
 	 	 	 	 <= GFF9BG
 	 	 	when 1000010111=> 
 	 	 	 	 <= GEE98C
 	 	 	when 1000011000=> 
 	 	 	 	 <= GDD762
 	 	 	when 1000011001=> 
 	 	 	 	 <= GBC538
 	 	 	when 1000011010=> 
 	 	 	 	 <= G9B30G
 	 	 	when 1000011011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000011100=> 
 	 	 	 	 <= GFFBC2
 	 	 	when 1000011101=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1000011110=> 
 	 	 	 	 <= G9B719
 	 	 	when 1000100000=> 
 	 	 	 	 <= GBC745
 	 	 	when 1000100001=> 
 	 	 	 	 <= G99E01
 	 	 	when 1000100010=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1000100011=> 
 	 	 	 	 <= GFF6B8
 	 	 	when 1000100100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000100101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000100110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000100111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000101000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000101001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000101010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000101011=> 
 	 	 	 	 <= G9B91D
 	 	 	when 1000101100=> 
 	 	 	 	 <= GEEG99
 	 	 	when 1000101101=> 
 	 	 	 	 <= GDE076
 	 	 	when 1000101110=> 
 	 	 	 	 <= G9B008
 	 	 	when 1000101111=> 
 	 	 	 	 <= GEEG98
 	 	 	when 1000110000=> 
 	 	 	 	 <= GEF29G
 	 	 	when 1000110001=> 
 	 	 	 	 <= GFFBC2
 	 	 	when 1000110010=> 
 	 	 	 	 <= G9B411
 	 	 	when 1000110011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000110100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000110101=> 
 	 	 	 	 <= G99D00
 	 	 	when 1000110110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000110111=> 
 	 	 	 	 <= G9B91E
 	 	 	when 1000111000=> 
 	 	 	 	 <= GCCC46
 	 	 	when 1000111001=> 
 	 	 	 	 <= GDDE70
 	 	 	when 1000111010=> 
 	 	 	 	 <= GEEG99
 	 	 	when 1000111011=> 
 	 	 	 	 <= GFFDC7
 	 	 	when 1000111100=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1000111101=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1000111110=> 
 	 	 	 	 <= G99G06
 	 	 	when 1001000000=> 
 	 	 	 	 <= GCD870
 	 	 	when 1001000001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001000010=> 
 	 	 	 	 <= GFF3B2
 	 	 	when 1001000011=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1001000100=> 
 	 	 	 	 <= G9B10B
 	 	 	when 1001000101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001000110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001000111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001001000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001001001=> 
 	 	 	 	 <= G99E01
 	 	 	when 1001001010=> 
 	 	 	 	 <= GCD55D
 	 	 	when 1001001011=> 
 	 	 	 	 <= GFF5B7
 	 	 	when 1001001100=> 
 	 	 	 	 <= GBC230
 	 	 	when 1001001101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001001110=> 
 	 	 	 	 <= G99D00
 	 	 	when 1001001111=> 
 	 	 	 	 <= GFF9BG
 	 	 	when 1001010000=> 
 	 	 	 	 <= G9B008
 	 	 	when 1001010001=> 
 	 	 	 	 <= GCC940
 	 	 	when 1001010010=> 
 	 	 	 	 <= GEEF97
 	 	 	when 1001010011=> 
 	 	 	 	 <= G99E02
 	 	 	when 1001010100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001010101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001010110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001010111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001011000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001011001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001011010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001011011=> 
 	 	 	 	 <= GCCC46
 	 	 	when 1001011100=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1001011101=> 
 	 	 	 	 <= GFF7BD
 	 	 	when 1001011110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001100000=> 
 	 	 	 	 <= GEF0C0
 	 	 	when 1001100001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001100010=> 
 	 	 	 	 <= GDDC6B
 	 	 	when 1001100011=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1001100100=> 
 	 	 	 	 <= GCCD47
 	 	 	when 1001100101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001100110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001100111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001101000=> 
 	 	 	 	 <= GBBC21
 	 	 	when 1001101001=> 
 	 	 	 	 <= GEF19F
 	 	 	when 1001101010=> 
 	 	 	 	 <= GDDE6G
 	 	 	when 1001101011=> 
 	 	 	 	 <= G99G06
 	 	 	when 1001101100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001101101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001101110=> 
 	 	 	 	 <= G9B411
 	 	 	when 1001101111=> 
 	 	 	 	 <= GFF3B3
 	 	 	when 1001110000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001110001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001110010=> 
 	 	 	 	 <= GDDE6G
 	 	 	when 1001110011=> 
 	 	 	 	 <= GDDD6E
 	 	 	when 1001110100=> 
 	 	 	 	 <= G99D00
 	 	 	when 1001110101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001110110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001110111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001111000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001111001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001111010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001111011=> 
 	 	 	 	 <= GCC941
 	 	 	when 1001111100=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1001111101=> 
 	 	 	 	 <= GDDG74
 	 	 	when 1001111110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010000000=> 
 	 	 	 	 <= GFGCG6
 	 	 	when 1010000001=> 
 	 	 	 	 <= G99G06
 	 	 	when 1010000010=> 
 	 	 	 	 <= G9BB20
 	 	 	when 1010000011=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1010000100=> 
 	 	 	 	 <= GFF3B2
 	 	 	when 1010000101=> 
 	 	 	 	 <= G9B615
 	 	 	when 1010000110=> 
 	 	 	 	 <= G99F03
 	 	 	when 1010000111=> 
 	 	 	 	 <= GDD863
 	 	 	when 1010001000=> 
 	 	 	 	 <= GFF4B4
 	 	 	when 1010001001=> 
 	 	 	 	 <= GBBG2B
 	 	 	when 1010001010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010001011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010001100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010001101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010001110=> 
 	 	 	 	 <= GBC840
 	 	 	when 1010001111=> 
 	 	 	 	 <= GDDG74
 	 	 	when 1010010000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010010001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010010010=> 
 	 	 	 	 <= G99F02
 	 	 	when 1010010011=> 
 	 	 	 	 <= GEEG98
 	 	 	when 1010010100=> 
 	 	 	 	 <= GCC83G
 	 	 	when 1010010101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010010110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010010111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010011000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010011001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010011010=> 
 	 	 	 	 <= G89D00
 	 	 	when 1010011011=> 
 	 	 	 	 <= GEEE94
 	 	 	when 1010011100=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 1010011101=> 
 	 	 	 	 <= GBBG2B
 	 	 	when 1010011110=> 
 	 	 	 	 <= G89D00
 	 	 	when 1010100001=> 
 	 	 	 	 <= GCD261
 	 	 	when 1010100010=> 
 	 	 	 	 <= G99D00
 	 	 	when 1010100011=> 
 	 	 	 	 <= GEEB8F
 	 	 	when 1010100100=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1010100101=> 
 	 	 	 	 <= GFFBC1
 	 	 	when 1010100110=> 
 	 	 	 	 <= GFF5B7
 	 	 	when 1010100111=> 
 	 	 	 	 <= GDDB68
 	 	 	when 1010101000=> 
 	 	 	 	 <= G99F04
 	 	 	when 1010101001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010101010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010101011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010101100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010101101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010101110=> 
 	 	 	 	 <= GDDE6F
 	 	 	when 1010101111=> 
 	 	 	 	 <= GCCC45
 	 	 	when 1010110000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010110001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010110010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010110011=> 
 	 	 	 	 <= G9B412
 	 	 	when 1010110100=> 
 	 	 	 	 <= GFF7BD
 	 	 	when 1010110101=> 
 	 	 	 	 <= G9B81C
 	 	 	when 1010110110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010110111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010111000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010111001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010111010=> 
 	 	 	 	 <= GBC537
 	 	 	when 1010111011=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1010111100=> 
 	 	 	 	 <= GEEG98
 	 	 	when 1010111101=> 
 	 	 	 	 <= G99D00
 	 	 	when 1010111110=> 
 	 	 	 	 <= GBC033
 	 	 	when 1011000001=> 
 	 	 	 	 <= GFG2EG
 	 	 	when 1011000010=> 
 	 	 	 	 <= G99F02
 	 	 	when 1011000011=> 
 	 	 	 	 <= G9B91F
 	 	 	when 1011000100=> 
 	 	 	 	 <= GFFGCF
 	 	 	when 1011000101=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1011000110=> 
 	 	 	 	 <= GDDG74
 	 	 	when 1011000111=> 
 	 	 	 	 <= G99D00
 	 	 	when 1011001000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011001001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011001010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011001011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011001100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011001101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011001110=> 
 	 	 	 	 <= GEF19E
 	 	 	when 1011001111=> 
 	 	 	 	 <= G9B616
 	 	 	when 1011010000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011010001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011010010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011010011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011010100=> 
 	 	 	 	 <= GBC230
 	 	 	when 1011010101=> 
 	 	 	 	 <= GFF3B3
 	 	 	when 1011010110=> 
 	 	 	 	 <= G99G06
 	 	 	when 1011010111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011011000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011011001=> 
 	 	 	 	 <= G9B30F
 	 	 	when 1011011010=> 
 	 	 	 	 <= GFF9C0
 	 	 	when 1011011011=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1011011100=> 
 	 	 	 	 <= GBBE26
 	 	 	when 1011011101=> 
 	 	 	 	 <= G89D00
 	 	 	when 1011011110=> 
 	 	 	 	 <= GEF3C8
 	 	 	when 1011100001=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1011100010=> 
 	 	 	 	 <= GCDB77
 	 	 	when 1011100011=> 
 	 	 	 	 <= G99D00
 	 	 	when 1011100100=> 
 	 	 	 	 <= GCD154
 	 	 	when 1011100101=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1011100110=> 
 	 	 	 	 <= GFFCC5
 	 	 	when 1011100111=> 
 	 	 	 	 <= G9B20E
 	 	 	when 1011101000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011101001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011101010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011101011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011101100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011101101=> 
 	 	 	 	 <= G99F04
 	 	 	when 1011101110=> 
 	 	 	 	 <= GFFBC3
 	 	 	when 1011101111=> 
 	 	 	 	 <= G89E00
 	 	 	when 1011110000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011110001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011110010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011110011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011110100=> 
 	 	 	 	 <= G89E00
 	 	 	when 1011110101=> 
 	 	 	 	 <= GCD55D
 	 	 	when 1011110110=> 
 	 	 	 	 <= GDE47G
 	 	 	when 1011110111=> 
 	 	 	 	 <= G99D00
 	 	 	when 1011111000=> 
 	 	 	 	 <= G9B109
 	 	 	when 1011111001=> 
 	 	 	 	 <= GEF19D
 	 	 	when 1011111010=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1011111011=> 
 	 	 	 	 <= GDD761
 	 	 	when 1011111100=> 
 	 	 	 	 <= G99D00
 	 	 	when 1011111101=> 
 	 	 	 	 <= GBC848
 	 	 	when 1011111110=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1100000010=> 
 	 	 	 	 <= GFGEGB
 	 	 	when 1100000011=> 
 	 	 	 	 <= GBBG30
 	 	 	when 1100000100=> 
 	 	 	 	 <= G99D00
 	 	 	when 1100000101=> 
 	 	 	 	 <= GDDG73
 	 	 	when 1100000110=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1100000111=> 
 	 	 	 	 <= GFF6B7
 	 	 	when 1100001000=> 
 	 	 	 	 <= G9B81C
 	 	 	when 1100001001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100001010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100001011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100001100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100001101=> 
 	 	 	 	 <= GBC02E
 	 	 	when 1100001110=> 
 	 	 	 	 <= GEE787
 	 	 	when 1100001111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100010000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100010001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100010010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100010011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100010100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100010101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100010110=> 
 	 	 	 	 <= GEE98C
 	 	 	when 1100010111=> 
 	 	 	 	 <= GEEC8G
 	 	 	when 1100011000=> 
 	 	 	 	 <= GFF7BB
 	 	 	when 1100011001=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1100011010=> 
 	 	 	 	 <= GDE37F
 	 	 	when 1100011011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100011100=> 
 	 	 	 	 <= G9B414
 	 	 	when 1100011101=> 
 	 	 	 	 <= GFG6FB
 	 	 	when 1100100011=> 
 	 	 	 	 <= GFG6F8
 	 	 	when 1100100100=> 
 	 	 	 	 <= G9B71B
 	 	 	when 1100100101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100100110=> 
 	 	 	 	 <= GDDC6D
 	 	 	when 1100100111=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1100101000=> 
 	 	 	 	 <= GFFFCC
 	 	 	when 1100101001=> 
 	 	 	 	 <= GCD358
 	 	 	when 1100101010=> 
 	 	 	 	 <= G99F03
 	 	 	when 1100101011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100101100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100101101=> 
 	 	 	 	 <= GCD55D
 	 	 	when 1100101110=> 
 	 	 	 	 <= GCD358
 	 	 	when 1100101111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100110000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100110001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100110010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100110011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100110100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100110101=> 
 	 	 	 	 <= G99F02
 	 	 	when 1100110110=> 
 	 	 	 	 <= GEE685
 	 	 	when 1100110111=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1100111000=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1100111001=> 
 	 	 	 	 <= GDDG73
 	 	 	when 1100111010=> 
 	 	 	 	 <= G99E01
 	 	 	when 1100111011=> 
 	 	 	 	 <= G9B008
 	 	 	when 1100111100=> 
 	 	 	 	 <= GEFCDD
 	 	 	when 1101000100=> 
 	 	 	 	 <= GFG3F0
 	 	 	when 1101000101=> 
 	 	 	 	 <= G9B91G
 	 	 	when 1101000110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1101000111=> 
 	 	 	 	 <= GBC83G
 	 	 	when 1101001000=> 
 	 	 	 	 <= GFFCC4
 	 	 	when 1101001001=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1101001010=> 
 	 	 	 	 <= GFFBC1
 	 	 	when 1101001011=> 
 	 	 	 	 <= GDD863
 	 	 	when 1101001100=> 
 	 	 	 	 <= GBC02D
 	 	 	when 1101001101=> 
 	 	 	 	 <= GFF3B1
 	 	 	when 1101001110=> 
 	 	 	 	 <= GCCF4F
 	 	 	when 1101001111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1101010000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1101010001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1101010010=> 
 	 	 	 	 <= G99D00
 	 	 	when 1101010011=> 
 	 	 	 	 <= G9B91E
 	 	 	when 1101010100=> 
 	 	 	 	 <= GCD65G
 	 	 	when 1101010101=> 
 	 	 	 	 <= GFF8BF
 	 	 	when 1101010110=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1101010111=> 
 	 	 	 	 <= GFFDC6
 	 	 	when 1101011000=> 
 	 	 	 	 <= GCCB44
 	 	 	when 1101011001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1101011010=> 
 	 	 	 	 <= G9B20E
 	 	 	when 1101011011=> 
 	 	 	 	 <= GEF9D7
 	 	 	when 1101100101=> 
 	 	 	 	 <= GFG8FG
 	 	 	when 1101100110=> 
 	 	 	 	 <= GBC846
 	 	 	when 1101100111=> 
 	 	 	 	 <= G99D00
 	 	 	when 1101101000=> 
 	 	 	 	 <= G9B10B
 	 	 	when 1101101001=> 
 	 	 	 	 <= GDD965
 	 	 	when 1101101010=> 
 	 	 	 	 <= GFFDC7
 	 	 	when 1101101011=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 1101101100=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1101101101=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1101101110=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1101101111=> 
 	 	 	 	 <= GFF2B0
 	 	 	when 1101110000=> 
 	 	 	 	 <= GEEE94
 	 	 	when 1101110001=> 
 	 	 	 	 <= GEF09C
 	 	 	when 1101110010=> 
 	 	 	 	 <= GFFEC8
 	 	 	when 1101110011=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1101110100=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1101110101=> 
 	 	 	 	 <= GFFEC9
 	 	 	when 1101110110=> 
 	 	 	 	 <= GDDC6B
 	 	 	when 1101110111=> 
 	 	 	 	 <= G9B20D
 	 	 	when 1101111000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1101111001=> 
 	 	 	 	 <= GBBG2G
 	 	 	when 1101111010=> 
 	 	 	 	 <= GFG3F0
 	 	 	when 1110000110=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1110000111=> 
 	 	 	 	 <= GDECB2
 	 	 	when 1110001000=> 
 	 	 	 	 <= G9B516
 	 	 	when 1110001001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1110001010=> 
 	 	 	 	 <= G99F04
 	 	 	when 1110001011=> 
 	 	 	 	 <= GBC73D
 	 	 	when 1110001100=> 
 	 	 	 	 <= GDE075
 	 	 	when 1110001101=> 
 	 	 	 	 <= GEF29G
 	 	 	when 1110001110=> 
 	 	 	 	 <= GFFFCC
 	 	 	when 1110001111=> 
 	 	 	 	 <= GGG0D1
 	 	 	when 1110010000=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1110010001=> 
 	 	 	 	 <= GFFFCD
 	 	 	when 1110010010=> 
 	 	 	 	 <= GFF3B1
 	 	 	when 1110010011=> 
 	 	 	 	 <= GDE178
 	 	 	when 1110010100=> 
 	 	 	 	 <= GBC840
 	 	 	when 1110010101=> 
 	 	 	 	 <= G99G05
 	 	 	when 1110010110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1110010111=> 
 	 	 	 	 <= G9B10C
 	 	 	when 1110011000=> 
 	 	 	 	 <= GDE188
 	 	 	when 1110011001=> 
 	 	 	 	 <= GFGEGD
 	 	 	when 1110101000=> 
 	 	 	 	 <= GFGEGB
 	 	 	when 1110101001=> 
 	 	 	 	 <= GDE99D
 	 	 	when 1110101010=> 
 	 	 	 	 <= GBC033
 	 	 	when 1110101011=> 
 	 	 	 	 <= G99D00
 	 	 	when 1110101100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1110101101=> 
 	 	 	 	 <= G89D00
 	 	 	when 1110101110=> 
 	 	 	 	 <= G99D00
 	 	 	when 1110101111=> 
 	 	 	 	 <= G99D00
 	 	 	when 1110110000=> 
 	 	 	 	 <= G99D00
 	 	 	when 1110110001=> 
 	 	 	 	 <= G89D00
 	 	 	when 1110110010=> 
 	 	 	 	 <= G89D00
 	 	 	when 1110110011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1110110100=> 
 	 	 	 	 <= G89D00
 	 	 	when 1110110101=> 
 	 	 	 	 <= G9BB22
 	 	 	when 1110110110=> 
 	 	 	 	 <= GDE188
 	 	 	when 1110110111=> 
 	 	 	 	 <= GFG9G1
 	 	 	when 1111001010=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1111001011=> 
 	 	 	 	 <= GFG6FB
 	 	 	when 1111001100=> 
 	 	 	 	 <= GDEEB8
 	 	 	when 1111001101=> 
 	 	 	 	 <= GCDB76
 	 	 	when 1111001110=> 
 	 	 	 	 <= GCCE54
 	 	 	when 1111001111=> 
 	 	 	 	 <= GBC643
 	 	 	when 1111010000=> 
 	 	 	 	 <= GBC642
 	 	 	when 1111010001=> 
 	 	 	 	 <= GBCD51
 	 	 	when 1111010010=> 
 	 	 	 	 <= GCD76F
 	 	 	when 1111010011=> 
 	 	 	 	 <= GDE99F
 	 	 	when 1111010100=> 
 	 	 	 	 <= GFG2EF
 	 	 	when 1111010101=> 
 	 	 	 	 <= GFGFGF 
 	 	 end case; 
     	 end if;  
     end process; 
 address <= row & col; 
 end;