library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ROM is
  port(
	  row : in std_logic_vector(4 downto 0);
	  col : in std_logic_vector(4 downto 0);
	  fruit_color : in std_logic_vector(5 downto 0);
	  clk : in std_logic;
	  color : out std_logic_vector(5 downto 0)
  );
end ROM;

architecture synth of ROM is 
signal address : std_logic_vector(9 downto 0);
begin
	process(clk) is
	begin
		if rising_edge(clk) then
			case address is 

 	 	 	when "0000000100010100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000000100010101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000000100010110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000000100010111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000001000010011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000001000010100" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0000001000010101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000001000010110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000001000010111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000001000011000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000001100010100" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0000001100010101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000001100010110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000001100010111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000001100011000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010000001101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000010000010011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000010000010100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000010000010101" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000010000010110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010000010111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010000011000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000010100001100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000010100001101" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000010100010100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000010100010101" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0000010100010110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000010100010111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000011000001011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0000011000001100" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000011000001101" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000011000010101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000011000010110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000011100001100" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000011100001101" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000100000001100" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0000100000001101" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000100000010010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0000100000010011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100000010100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100000010101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000100000101111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000100100010010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0000100100010011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100100010100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100100010101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100100101101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0000100100101110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0000100100101111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0000100100110000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0000100100110001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0000101000010001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101000010010" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000101000010011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101000010100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101000010101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101000010110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000101000100010" => 
 	 	 	 	 color <= "101011";
 	 	 	when "0000101000100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0000101000101011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000101000101100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0000101000101101" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000101000101110" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000101000101111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0000101000110000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000101000110001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0000101000110010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0000101100010001" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0000101100010010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000101100010011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101100010100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101100010101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101100010110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000101100100010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0000101100101011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0000101100101100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000101100101101" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0000101100101110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000101100101111" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0000101100110000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000101100110001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000101100110010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0000101100110011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000110000010001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000110000010010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110000010011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110000010100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110000010101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000110000100010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000110000100011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0000110000101010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000110000101011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0000110000101100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0000110000101101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000110000101110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000110000101111" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0000110000110000" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0000110000110001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000110000110010" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000110000110011" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0000110100100010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0000110100100011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0000110100101010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000110100101011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000110100101100" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0000110100101101" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0000110100101110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000110100101111" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000110100110000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000110100110001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000110100110010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000110100110011" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0000111000100010" => 
 	 	 	 	 color <= "101011";
 	 	 	when "0000111000100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0000111000101010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000111000101011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0000111000101100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000111000101101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000111000101110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000111000101111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000111000110000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000111000110001" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000111000110010" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000111000110011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0000111100100010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0000111100100011" => 
 	 	 	 	 color <= "101011";
 	 	 	when "0000111100101011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0000111100101100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000111100101101" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0000111100101110" => 
 	 	 	 	 color <= "110100";
 	 	 	when "0000111100101111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000111100110000" => 
 	 	 	 	 color <= "110000";
 	 	 	when "0000111100110001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0000111100110010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001000000100010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001000000100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001000000101011" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001000000101100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001000000101101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001000000101110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001000000101111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001000000110000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001000000110001" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0001000000110010" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0001000100100010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001000100100011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001000100101101" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0001000100101110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001000100101111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001000100110000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001000100110001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001001000010011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001001000100010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001001000100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001001100010010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001100010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001001100010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001001100010101" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0001001100011001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001001100011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001001100011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001001100011100" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001001100100010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001001100100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001010000010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001010000010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001010000010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001010000010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001010000010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001010000010111" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0001010000011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001010000011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001010000011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001010000011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001010000011101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0001010000011110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0001010000011111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001010000100010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0001010000100011" => 
 	 	 	 	 color <= "011010";
 	 	 	when "0001010100010001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001010100010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001010100010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001010100010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001010100010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001010100010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001010100010111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001010100011000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001010100011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001010100011010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001010100011011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001010100011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001010100011101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001010100011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001010100011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001010100100010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001010100100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001011000010010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001011000010011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001011000010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001011000010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001011000010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001011000010111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001011000011000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001011000011001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0001011000011010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001011000011011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001011000011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001011000011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001011000011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001011000011111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001011000100011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001011100010001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001011100010010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001011100010011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001011100010100" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0001011100010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001011100010110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001011100011000" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0001011100011001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001011100011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001011100011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001011100011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001011100011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001011100100010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0001011100100011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0001100000010000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100000010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001100000010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001100000010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001100000010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001100000010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001100000010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001100000010111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001100000011000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001100000011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001100000011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001100000011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001100000011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001100000011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001100000011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001100000011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0001100000100010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001100000100011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001100100010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001100100010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001100100010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001100100010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001100100010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001100100010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001100100010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001100100010111" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0001100100011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001100100011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001100100011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001100100011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001100100011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001100100011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001100100011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001100100100010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0001100100100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001100100100110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001101000010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001101000010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001101000010010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0001101000010011" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0001101000010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001101000010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001101000010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001101000010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001101000011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001101000011001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001101000011010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001101000011011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001101000011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001101000011101" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0001101000011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001101000100010" => 
 	 	 	 	 color <= "111011";
 	 	 	when "0001101000100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001101000100101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001101000100110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001101000100111" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001101100010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001101100010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001101100010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001101100010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001101100010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001101100010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001101100010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001101100010111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0001101100011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001101100011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001101100011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001101100011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001101100011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001101100011101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001101100100010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001101100100011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001101100100101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001101100100110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001101100100111" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001110000010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001110000010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001110000010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001110000010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001110000010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001110000010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001110000010111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110000011000" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0001110000011001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001110000011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001110000011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001110000011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001110000011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001110000100010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0001110000100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001110000100101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001110100000011" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0001110100000100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001110100000101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001110100000110" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0001110100010001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001110100010010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0001110100010011" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0001110100010100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001110100010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001110100010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001110100010111" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0001110100011000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001110100011001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0001110100011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001110100011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001110100011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001110100011101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001110100100010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001110100100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001110100100101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001110100100110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001110100100111" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001111000000010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001111000000011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001111000000100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001111000000101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001111000000110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001111000000111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001111000010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001111000010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001111000010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001111000010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001111000010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001111000010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001111000010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001111000010111" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001111000011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001111000011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001111000011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001111000011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001111000011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001111000011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001111000100010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0001111000100011" => 
 	 	 	 	 color <= "101011";
 	 	 	when "0001111000100110" => 
 	 	 	 	 color <= "011010";
 	 	 	when "0001111000100111" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001111100000001" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0001111100000010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001111100000011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001111100000100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001111100000101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001111100000110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0001111100000111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001111100001000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0001111100001111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001111100010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001111100010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001111100010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001111100010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001111100010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001111100010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001111100010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0001111100010111" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0001111100011000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001111100011001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001111100011010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001111100011011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0001111100011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001111100011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0001111100100101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0001111100100110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010000000000001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010000000000010" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0010000000000011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010000000000100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010000000000101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010000000000110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010000000000111" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0010000000001000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010000000010000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010000000010001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010000000010100" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010000000010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010000000010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010000000010111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000000011011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0010000000011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010000000011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010000000100010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010000000100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010000000100110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010000000100111" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010000100000001" => 
 	 	 	 	 color <= "111101";
 	 	 	when "0010000100000010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010000100000011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010000100000100" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000100000101" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000100000110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010000100000111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010000100001000" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010000100010000" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010000100010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010000100010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010000100010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010000100010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010000100010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010000100010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010000100010111" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010000100011001" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0010000100011010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0010000100011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010000100011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010000100011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010000100011110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0010000100100010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010000100100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010000100100101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010000100100110" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010000100100111" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010001000000001" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010001000000010" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010001000000011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010001000000100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010001000000101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010001000000110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010001000000111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010001000001000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010001000001111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001000010000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010001000010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010001000010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010001000010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010001000010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010001000010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010001000010110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010001000011000" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0010001000011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010001000011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010001000011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010001000011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010001000011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010001000011110" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0010001000100010" => 
 	 	 	 	 color <= "101011";
 	 	 	when "0010001000100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010001000100101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010001000100110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010001000100111" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010001100000001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010001100000010" => 
 	 	 	 	 color <= "111101";
 	 	 	when "0010001100000011" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0010001100000100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010001100000101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010001100000110" => 
 	 	 	 	 color <= "111000";
 	 	 	when "0010001100000111" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010001100001000" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010001100010000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001100010001" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010001100010010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010001100010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010001100010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010001100010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010001100010110" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010001100010111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0010001100011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010001100011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010001100011010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0010001100011011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0010001100011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010001100011101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0010001100100010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010001100100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010001100100110" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010010000000010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0010010000000011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010010000000100" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010010000000101" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010010000000110" => 
 	 	 	 	 color <= "111101";
 	 	 	when "0010010000000111" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0010010000010001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010010000010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010000010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010000010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010000010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010000010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010000010111" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0010010000011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010010000011001" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0010010000011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010010000011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010010000011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010010000011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010010000011110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0010010000100010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010010000100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010010000100101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010010000100110" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010010000100111" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010010100000100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010010100000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010010100010000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010010100010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010100010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010100010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010100010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010100010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010100010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010010100010111" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010010100011000" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010010100011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010010100011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010010100011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010010100011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010010100011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010010100011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010010100100010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010010100100101" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010011000010000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010011000010001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010011000010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010011000010011" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010011000010100" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0010011000010101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010011000011001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0010011000011010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0010011000011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010011000011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010011000011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010011000011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010011000011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0010011000100010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010011000100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010011100010001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010011100010010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010011100010110" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010011100010111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010011100011000" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010011100011001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0010011100011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010011100011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010011100011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010011100011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010011100011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010011100011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0010100000010001" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010100000010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100000010011" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0010100000010100" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010100000010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100000010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100000010111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100000011000" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010100000011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010100000011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010100000011011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0010100000011100" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0010100000011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010100000011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010100000011111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0010100000100010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010100000100011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010100100010001" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010100100010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100100010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100100010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100100010101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100100010110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100100010111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010100100011000" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0010100100011001" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010100100011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010100100011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010100100011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010100100011101" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010100100011110" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010100100011111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0010100100100010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010100100101101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0010101000010001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010101000010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010101000010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010101000010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010101000010101" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0010101000010110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010101000011010" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010101000011011" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010101000011100" => 
 	 	 	 	 color <= "101101";
 	 	 	when "0010101000011101" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0010101000011110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0010101000100010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010101000100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010101000101100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010101000101101" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010101000101110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0010101100010010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010101100010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010101100010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010101100100011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010101100101011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010101100101100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010101100101101" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010101100101110" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0010110000010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010110000010100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010110000100010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010110000100011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010110000101011" => 
 	 	 	 	 color <= "110001";
 	 	 	when "0010110000101100" => 
 	 	 	 	 color <= "100001";
 	 	 	when "0010110000101101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010110000101110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0010110000101111" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0010110100100010" => 
 	 	 	 	 color <= "111011";
 	 	 	when "0010110100100011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0010110100101010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010110100101011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010110100101100" => 
 	 	 	 	 color <= "100001";
 	 	 	when "0010110100101101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010110100101110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0010110100101111" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0010111000100010" => 
 	 	 	 	 color <= "011010";
 	 	 	when "0010111000100011" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010111000101001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010111000101010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010111000101011" => 
 	 	 	 	 color <= "100001";
 	 	 	when "0010111000101100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010111000101101" => 
 	 	 	 	 color <= "110001";
 	 	 	when "0010111000101110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010111000101111" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0010111100101001" => 
 	 	 	 	 color <= "100001";
 	 	 	when "0010111100101010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010111100101011" => 
 	 	 	 	 color <= "110001";
 	 	 	when "0010111100101100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010111100101101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010111100101110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010111100101111" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011000000101000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0011000000101001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011000000101010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011000000101011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011000000101100" => 
 	 	 	 	 color <= "110001";
 	 	 	when "0011000000101101" => 
 	 	 	 	 color <= "110001";
 	 	 	when "0011000000101110" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0011000000101111" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0011000100100010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011000100100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011000100101000" => 
 	 	 	 	 color <= "110001";
 	 	 	when "0011000100101001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011000100101010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011000100101011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011000100101100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011000100101101" => 
 	 	 	 	 color <= "110001";
 	 	 	when "0011000100101110" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011000100101111" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0011001000001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011001000001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011001000001111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0011001000100111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011001000101000" => 
 	 	 	 	 color <= "100001";
 	 	 	when "0011001000101001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011001000101010" => 
 	 	 	 	 color <= "110001";
 	 	 	when "0011001000101011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011001000101100" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011001000101101" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0011001000101110" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0011001100001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011001100001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011001100001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011001100001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011001100100010" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011001100100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011001100100111" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011001100101000" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011001100101001" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011001100101010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011001100101011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011001100101100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0011001100101101" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011001100101110" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0011010000001001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0011010000001010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0011010000001011" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011010000001100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0011010000001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011010000001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011010000001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011010000010000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0011010000100010" => 
 	 	 	 	 color <= "010101";
 	 	 	when "0011010000100011" => 
 	 	 	 	 color <= "101010";
 	 	 	when "0011010000100110" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0011010000100111" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010000101000" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0011010000101001" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0011010000101010" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010000101011" => 
 	 	 	 	 color <= "111110";
 	 	 	when "0011010000101100" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0011010000101101" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0011010100001010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0011010100001011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0011010100001100" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0011010100001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011010100001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011010100001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011010100010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011010100010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011010100100010" => 
 	 	 	 	 color <= "010001";
 	 	 	when "0011010100100111" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0011010100101000" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0011010100101001" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0011010100101010" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0011010100101011" => 
 	 	 	 	 color <= "000100";
 	 	 	when "0011011000001010" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0011011000001011" => 
 	 	 	 	 color <= "011001";
 	 	 	when "0011011000001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011000001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011000001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011000001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011000010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011000010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011000010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011100001001" => 
 	 	 	 	 color <= "010100";
 	 	 	when "0011011100001010" => 
 	 	 	 	 color <= "101001";
 	 	 	when "0011011100001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011100001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011100001101" => 
 	 	 	 	 color <= "000110";
 	 	 	when "0011011100001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011100001111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0011011100010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011100010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011100010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011100010011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0011100000001010" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0011100000001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100000001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100000001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100000001110" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0011100000001111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0011100000010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100000010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100000010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100000010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100100001011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0011100100001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100100001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100100001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100100001111" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0011100100010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100100010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100100010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100100010011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0011101000001011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0011101000001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011101000001101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0011101000001110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0011101000001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011101000010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011101000010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011101000010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011101100010000" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0011101100010001" => 
 	 	 	 	 color <= "000001"; 
 	 	 end case; 
     	 end if;  
     end process; 
 address <= row & col; 
 end;