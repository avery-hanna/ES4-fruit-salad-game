library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity WATERMELONROM is
  port(
	  row : in std_logic_vector(4 downto 0);
	  col : in std_logic_vector(4 downto 0);
	  fruit_color : in std_logic_vector(5 downto 0);
	  clk : in std_logic;
	  color : out std_logic_vector(5 downto 0)
  );
end WATERMELONROM;

architecture synth of WATERMELONROM is 
signal address : std_logic_vector(9 downto 0);
begin
	process(clk) is
	begin
		if rising_edge(clk) then
			case address is 

 	 	 	when 0000001100=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000001101=> 
 	 	 	 	 <= GDGEGE
 	 	 	when 0000001110=> 
 	 	 	 	 <= F4G0FB
 	 	 	when 0000001111=> 
 	 	 	 	 <= EBFBF2
 	 	 	when 0000010000=> 
 	 	 	 	 <= EEFDF4
 	 	 	when 0000010001=> 
 	 	 	 	 <= G3G8G6
 	 	 	when 0000010010=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000101001=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000101010=> 
 	 	 	 	 <= D8F1E4
 	 	 	when 0000101011=> 
 	 	 	 	 <= 6FBG8G
 	 	 	when 0000101100=> 
 	 	 	 	 <= 288959
 	 	 	when 0000101101=> 
 	 	 	 	 <= 01733B
 	 	 	when 0000101110=> 
 	 	 	 	 <= 007339
 	 	 	when 0000101111=> 
 	 	 	 	 <= 00723B
 	 	 	when 0000110000=> 
 	 	 	 	 <= 00733B
 	 	 	when 0000110001=> 
 	 	 	 	 <= 00723B
 	 	 	when 0000110010=> 
 	 	 	 	 <= 0F7B45
 	 	 	when 0000110011=> 
 	 	 	 	 <= 4B9C73
 	 	 	when 0000110100=> 
 	 	 	 	 <= 9CD8C1
 	 	 	when 0000110101=> 
 	 	 	 	 <= G3G8G5
 	 	 	when 0001000111=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0001001000=> 
 	 	 	 	 <= C2E5D4
 	 	 	when 0001001001=> 
 	 	 	 	 <= 2C8B5C
 	 	 	when 0001001010=> 
 	 	 	 	 <= 00733B
 	 	 	when 0001001011=> 
 	 	 	 	 <= 00733B
 	 	 	when 0001001100=> 
 	 	 	 	 <= 05753E
 	 	 	when 0001001101=> 
 	 	 	 	 <= 32885C
 	 	 	when 0001001110=> 
 	 	 	 	 <= 549771
 	 	 	when 0001001111=> 
 	 	 	 	 <= 609D79
 	 	 	when 0001010000=> 
 	 	 	 	 <= 599974
 	 	 	when 0001010001=> 
 	 	 	 	 <= 3D8E61
 	 	 	when 0001010010=> 
 	 	 	 	 <= 0E7842
 	 	 	when 0001010011=> 
 	 	 	 	 <= 00733B
 	 	 	when 0001010100=> 
 	 	 	 	 <= 00733B
 	 	 	when 0001010101=> 
 	 	 	 	 <= 077740
 	 	 	when 0001010110=> 
 	 	 	 	 <= 72C192
 	 	 	when 0001010111=> 
 	 	 	 	 <= G0G6G3
 	 	 	when 0001100110=> 
 	 	 	 	 <= FCG4G0
 	 	 	when 0001100111=> 
 	 	 	 	 <= 489B71
 	 	 	when 0001101000=> 
 	 	 	 	 <= 00723B
 	 	 	when 0001101001=> 
 	 	 	 	 <= 01733C
 	 	 	when 0001101010=> 
 	 	 	 	 <= 549771
 	 	 	when 0001101011=> 
 	 	 	 	 <= C8C8B9
 	 	 	when 0001101100=> 
 	 	 	 	 <= FGBFBF
 	 	 	when 0001101101=> 
 	 	 	 	 <= FD9595
 	 	 	when 0001101110=> 
 	 	 	 	 <= F88484
 	 	 	when 0001101111=> 
 	 	 	 	 <= F77G7G
 	 	 	when 0001110000=> 
 	 	 	 	 <= F78282
 	 	 	when 0001110001=> 
 	 	 	 	 <= FC9090
 	 	 	when 0001110010=> 
 	 	 	 	 <= G1B8B8
 	 	 	when 0001110011=> 
 	 	 	 	 <= DCC8BE
 	 	 	when 0001110100=> 
 	 	 	 	 <= 72B485
 	 	 	when 0001110101=> 
 	 	 	 	 <= 0D7842
 	 	 	when 0001110110=> 
 	 	 	 	 <= 00733B
 	 	 	when 0001110111=> 
 	 	 	 	 <= 107D46
 	 	 	when 0001111000=> 
 	 	 	 	 <= BDE1CG
 	 	 	when 0001111001=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0010000101=> 
 	 	 	 	 <= E2F6ED
 	 	 	when 0010000110=> 
 	 	 	 	 <= 177G4C
 	 	 	when 0010000111=> 
 	 	 	 	 <= 00733B
 	 	 	when 0010001000=> 
 	 	 	 	 <= 449066
 	 	 	when 0010001001=> 
 	 	 	 	 <= E7CCC3
 	 	 	when 0010001010=> 
 	 	 	 	 <= F98B8B
 	 	 	when 0010001011=> 
 	 	 	 	 <= F16969
 	 	 	when 0010001100=> 
 	 	 	 	 <= 7C3B3B
 	 	 	when 0010001101=> 
 	 	 	 	 <= CD5858
 	 	 	when 0010001110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0010001111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0010010000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0010010001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0010010010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0010010011=> 
 	 	 	 	 <= F1696B
 	 	 	when 0010010100=> 
 	 	 	 	 <= F67D7D
 	 	 	when 0010010101=> 
 	 	 	 	 <= F8C3C0
 	 	 	when 0010010110=> 
 	 	 	 	 <= 70B383
 	 	 	when 0010010111=> 
 	 	 	 	 <= 01733C
 	 	 	when 0010011000=> 
 	 	 	 	 <= 007239
 	 	 	when 0010011001=> 
 	 	 	 	 <= 74C293
 	 	 	when 0010011010=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0010100100=> 
 	 	 	 	 <= E2F6ED
 	 	 	when 0010100101=> 
 	 	 	 	 <= 0D7943
 	 	 	when 0010100110=> 
 	 	 	 	 <= 01733C
 	 	 	when 0010100111=> 
 	 	 	 	 <= 8GBF96
 	 	 	when 0010101000=> 
 	 	 	 	 <= FE9C9C
 	 	 	when 0010101001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0010101010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0010101011=> 
 	 	 	 	 <= F16969
 	 	 	when 0010101100=> 
 	 	 	 	 <= 572829
 	 	 	when 0010101101=> 
 	 	 	 	 <= 5F2D2D
 	 	 	when 0010101110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0010101111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0010110000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0010110001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0010110010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0010110011=> 
 	 	 	 	 <= 442020
 	 	 	when 0010110100=> 
 	 	 	 	 <= 5F2D2D
 	 	 	when 0010110101=> 
 	 	 	 	 <= F16969
 	 	 	when 0010110110=> 
 	 	 	 	 <= F88585
 	 	 	when 0010110111=> 
 	 	 	 	 <= D1CCBF
 	 	 	when 0010111000=> 
 	 	 	 	 <= 127B45
 	 	 	when 0010111001=> 
 	 	 	 	 <= 00723B
 	 	 	when 0010111010=> 
 	 	 	 	 <= 66BC89
 	 	 	when 0010111011=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0011000011=> 
 	 	 	 	 <= FBG3FG
 	 	 	when 0011000100=> 
 	 	 	 	 <= 167G4C
 	 	 	when 0011000101=> 
 	 	 	 	 <= 02733C
 	 	 	when 0011000110=> 
 	 	 	 	 <= BCC7B4
 	 	 	when 0011000111=> 
 	 	 	 	 <= F78282
 	 	 	when 0011001000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011001001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011001010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011001011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011001100=> 
 	 	 	 	 <= F16969
 	 	 	when 0011001101=> 
 	 	 	 	 <= F2696B
 	 	 	when 0011001110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011001111=> 
 	 	 	 	 <= DE6060
 	 	 	when 0011010000=> 
 	 	 	 	 <= F1696B
 	 	 	when 0011010001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011010010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011010011=> 
 	 	 	 	 <= C55454
 	 	 	when 0011010100=> 
 	 	 	 	 <= 622F2F
 	 	 	when 0011010101=> 
 	 	 	 	 <= EF6868
 	 	 	when 0011010110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011010111=> 
 	 	 	 	 <= F47272
 	 	 	when 0011011000=> 
 	 	 	 	 <= E8CCC4
 	 	 	when 0011011001=> 
 	 	 	 	 <= 167D48
 	 	 	when 0011011010=> 
 	 	 	 	 <= 007239
 	 	 	when 0011011011=> 
 	 	 	 	 <= 8CCGB5
 	 	 	when 0011011100=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0011100010=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0011100011=> 
 	 	 	 	 <= 469970
 	 	 	when 0011100100=> 
 	 	 	 	 <= 007239
 	 	 	when 0011100101=> 
 	 	 	 	 <= 96C099
 	 	 	when 0011100110=> 
 	 	 	 	 <= F78181
 	 	 	when 0011100111=> 
 	 	 	 	 <= F2696B
 	 	 	when 0011101000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011101001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011101010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011101011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011101100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011101101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011101110=> 
 	 	 	 	 <= DG6161
 	 	 	when 0011101111=> 
 	 	 	 	 <= 070303
 	 	 	when 0011110000=> 
 	 	 	 	 <= 4E2424
 	 	 	when 0011110001=> 
 	 	 	 	 <= F26969
 	 	 	when 0011110010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011110011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011110100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011110101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011110110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011110111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0011111000=> 
 	 	 	 	 <= F37070
 	 	 	when 0011111001=> 
 	 	 	 	 <= DFCDC2
 	 	 	when 0011111010=> 
 	 	 	 	 <= 06753F
 	 	 	when 0011111011=> 
 	 	 	 	 <= 02743C
 	 	 	when 0011111100=> 
 	 	 	 	 <= E0F5EB
 	 	 	when 0100000010=> 
 	 	 	 	 <= C0E4D2
 	 	 	when 0100000011=> 
 	 	 	 	 <= 007239
 	 	 	when 0100000100=> 
 	 	 	 	 <= 4E946D
 	 	 	when 0100000101=> 
 	 	 	 	 <= FD9696
 	 	 	when 0100000110=> 
 	 	 	 	 <= F16969
 	 	 	when 0100000111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100001000=> 
 	 	 	 	 <= 873G3G
 	 	 	when 0100001001=> 
 	 	 	 	 <= 994747
 	 	 	when 0100001010=> 
 	 	 	 	 <= F16969
 	 	 	when 0100001011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100001100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100001101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100001110=> 
 	 	 	 	 <= F2696B
 	 	 	when 0100001111=> 
 	 	 	 	 <= E26262
 	 	 	when 0100010000=> 
 	 	 	 	 <= CD5858
 	 	 	when 0100010001=> 
 	 	 	 	 <= F26B69
 	 	 	when 0100010010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100010011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100010100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100010101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100010110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100010111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100011000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100011001=> 
 	 	 	 	 <= F67B7B
 	 	 	when 0100011010=> 
 	 	 	 	 <= 94C098
 	 	 	when 0100011011=> 
 	 	 	 	 <= 00733B
 	 	 	when 0100011100=> 
 	 	 	 	 <= 328F61
 	 	 	when 0100011101=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0100100001=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0100100010=> 
 	 	 	 	 <= 278858
 	 	 	when 0100100011=> 
 	 	 	 	 <= 05753E
 	 	 	when 0100100100=> 
 	 	 	 	 <= EEC9C3
 	 	 	when 0100100101=> 
 	 	 	 	 <= F16B6B
 	 	 	when 0100100110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100100111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100101000=> 
 	 	 	 	 <= 763737
 	 	 	when 0100101001=> 
 	 	 	 	 <= 170B0B
 	 	 	when 0100101010=> 
 	 	 	 	 <= B44E4E
 	 	 	when 0100101011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100101100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100101101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100101110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100101111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100110000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100110001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100110010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100110011=> 
 	 	 	 	 <= F16969
 	 	 	when 0100110100=> 
 	 	 	 	 <= 8B4040
 	 	 	when 0100110101=> 
 	 	 	 	 <= 6D3233
 	 	 	when 0100110110=> 
 	 	 	 	 <= EF6868
 	 	 	when 0100110111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100111000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0100111001=> 
 	 	 	 	 <= F2696B
 	 	 	when 0100111010=> 
 	 	 	 	 <= FGB2B2
 	 	 	when 0100111011=> 
 	 	 	 	 <= 2C8556
 	 	 	when 0100111100=> 
 	 	 	 	 <= 007239
 	 	 	when 0100111101=> 
 	 	 	 	 <= C6E7D7
 	 	 	when 0101000001=> 
 	 	 	 	 <= D2EEE0
 	 	 	when 0101000010=> 
 	 	 	 	 <= 00733B
 	 	 	when 0101000011=> 
 	 	 	 	 <= 649F7D
 	 	 	when 0101000100=> 
 	 	 	 	 <= F88383
 	 	 	when 0101000101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101000110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101000111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101001000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101001001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101001010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101001011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101001100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101001101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101001110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101001111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101010000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101010001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101010010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101010011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101010100=> 
 	 	 	 	 <= C85656
 	 	 	when 0101010101=> 
 	 	 	 	 <= 4D2323
 	 	 	when 0101010110=> 
 	 	 	 	 <= DE6060
 	 	 	when 0101010111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101011000=> 
 	 	 	 	 <= E36363
 	 	 	when 0101011001=> 
 	 	 	 	 <= 5E2C2C
 	 	 	when 0101011010=> 
 	 	 	 	 <= D35F5G
 	 	 	when 0101011011=> 
 	 	 	 	 <= BCC6B4
 	 	 	when 0101011100=> 
 	 	 	 	 <= 00733B
 	 	 	when 0101011101=> 
 	 	 	 	 <= 45986G
 	 	 	when 0101011110=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0101100001=> 
 	 	 	 	 <= 67BC89
 	 	 	when 0101100010=> 
 	 	 	 	 <= 00733B
 	 	 	when 0101100011=> 
 	 	 	 	 <= D8C8BE
 	 	 	when 0101100100=> 
 	 	 	 	 <= F1696B
 	 	 	when 0101100101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101100110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101100111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101101000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101101001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101101010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101101011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101101100=> 
 	 	 	 	 <= F1696B
 	 	 	when 0101101101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101101110=> 
 	 	 	 	 <= F2696B
 	 	 	when 0101101111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101110000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101110001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101110010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101110011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101110100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101110101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101110110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101110111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0101111000=> 
 	 	 	 	 <= EC6666
 	 	 	when 0101111001=> 
 	 	 	 	 <= 472121
 	 	 	when 0101111010=> 
 	 	 	 	 <= 2D1415
 	 	 	when 0101111011=> 
 	 	 	 	 <= FGBCBC
 	 	 	when 0101111100=> 
 	 	 	 	 <= 0F7943
 	 	 	when 0101111101=> 
 	 	 	 	 <= 01733C
 	 	 	when 0101111110=> 
 	 	 	 	 <= G2G7G5
 	 	 	when 0110000000=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0110000001=> 
 	 	 	 	 <= 208453
 	 	 	when 0110000010=> 
 	 	 	 	 <= 117B45
 	 	 	when 0110000011=> 
 	 	 	 	 <= G0B7B7
 	 	 	when 0110000100=> 
 	 	 	 	 <= DG6161
 	 	 	when 0110000101=> 
 	 	 	 	 <= DC5G5G
 	 	 	when 0110000110=> 
 	 	 	 	 <= F26B69
 	 	 	when 0110000111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110001000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110001001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110001010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110001011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110001100=> 
 	 	 	 	 <= C65555
 	 	 	when 0110001101=> 
 	 	 	 	 <= 040202
 	 	 	when 0110001110=> 
 	 	 	 	 <= 843F3F
 	 	 	when 0110001111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110010000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110010001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110010010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110010011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110010100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110010101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110010110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110010111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110011000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110011001=> 
 	 	 	 	 <= F16B6B
 	 	 	when 0110011010=> 
 	 	 	 	 <= F1696B
 	 	 	when 0110011011=> 
 	 	 	 	 <= F88585
 	 	 	when 0110011100=> 
 	 	 	 	 <= 589873
 	 	 	when 0110011101=> 
 	 	 	 	 <= 007239
 	 	 	when 0110011110=> 
 	 	 	 	 <= C2E4D3
 	 	 	when 0110100000=> 
 	 	 	 	 <= G8GCGB
 	 	 	when 0110100001=> 
 	 	 	 	 <= 00733B
 	 	 	when 0110100010=> 
 	 	 	 	 <= 489269
 	 	 	when 0110100011=> 
 	 	 	 	 <= FB8C8C
 	 	 	when 0110100100=> 
 	 	 	 	 <= 713535
 	 	 	when 0110100101=> 
 	 	 	 	 <= 050202
 	 	 	when 0110100110=> 
 	 	 	 	 <= E86565
 	 	 	when 0110100111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110101000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110101001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110101010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110101011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110101100=> 
 	 	 	 	 <= F2696B
 	 	 	when 0110101101=> 
 	 	 	 	 <= C05252
 	 	 	when 0110101110=> 
 	 	 	 	 <= C25353
 	 	 	when 0110101111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110110000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110110001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110110010=> 
 	 	 	 	 <= C05252
 	 	 	when 0110110011=> 
 	 	 	 	 <= D45D5D
 	 	 	when 0110110100=> 
 	 	 	 	 <= F1696B
 	 	 	when 0110110101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110110110=> 
 	 	 	 	 <= F1696B
 	 	 	when 0110110111=> 
 	 	 	 	 <= 773838
 	 	 	when 0110111000=> 
 	 	 	 	 <= C75556
 	 	 	when 0110111001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110111010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0110111011=> 
 	 	 	 	 <= F26D6D
 	 	 	when 0110111100=> 
 	 	 	 	 <= 92C199
 	 	 	when 0110111101=> 
 	 	 	 	 <= 00733B
 	 	 	when 0110111110=> 
 	 	 	 	 <= 7GC89D
 	 	 	when 0111000000=> 
 	 	 	 	 <= EEFDF4
 	 	 	when 0111000001=> 
 	 	 	 	 <= 00733B
 	 	 	when 0111000010=> 
 	 	 	 	 <= 6EB281
 	 	 	when 0111000011=> 
 	 	 	 	 <= F57979
 	 	 	when 0111000100=> 
 	 	 	 	 <= F2696B
 	 	 	when 0111000101=> 
 	 	 	 	 <= F1696B
 	 	 	when 0111000110=> 
 	 	 	 	 <= F2696B
 	 	 	when 0111000111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111001000=> 
 	 	 	 	 <= F1696B
 	 	 	when 0111001001=> 
 	 	 	 	 <= F16B69
 	 	 	when 0111001010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111001011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111001100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111001101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111001110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111001111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111010000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111010001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111010010=> 
 	 	 	 	 <= 542727
 	 	 	when 0111010011=> 
 	 	 	 	 <= 150B0B
 	 	 	when 0111010100=> 
 	 	 	 	 <= EF6868
 	 	 	when 0111010101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111010110=> 
 	 	 	 	 <= F1696B
 	 	 	when 0111010111=> 
 	 	 	 	 <= 472121
 	 	 	when 0111011000=> 
 	 	 	 	 <= 090404
 	 	 	when 0111011001=> 
 	 	 	 	 <= EG6868
 	 	 	when 0111011010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111011011=> 
 	 	 	 	 <= F26969
 	 	 	when 0111011100=> 
 	 	 	 	 <= C3C6B6
 	 	 	when 0111011101=> 
 	 	 	 	 <= 00733B
 	 	 	when 0111011110=> 
 	 	 	 	 <= 5FB683
 	 	 	when 0111100000=> 
 	 	 	 	 <= DGF4EB
 	 	 	when 0111100001=> 
 	 	 	 	 <= 007239
 	 	 	when 0111100010=> 
 	 	 	 	 <= 7EB98D
 	 	 	when 0111100011=> 
 	 	 	 	 <= F37171
 	 	 	when 0111100100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111100101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111100110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111100111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111101000=> 
 	 	 	 	 <= 863F3G
 	 	 	when 0111101001=> 
 	 	 	 	 <= 160B0B
 	 	 	when 0111101010=> 
 	 	 	 	 <= BG5252
 	 	 	when 0111101011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111101100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111101101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111101110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111101111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111110000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111110001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111110010=> 
 	 	 	 	 <= F1696B
 	 	 	when 0111110011=> 
 	 	 	 	 <= F1696B
 	 	 	when 0111110100=> 
 	 	 	 	 <= F1696B
 	 	 	when 0111110101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111110110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111110111=> 
 	 	 	 	 <= F1696B
 	 	 	when 0111111000=> 
 	 	 	 	 <= F1696B
 	 	 	when 0111111001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111111010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 0111111011=> 
 	 	 	 	 <= F2696B
 	 	 	when 0111111100=> 
 	 	 	 	 <= CFC4B7
 	 	 	when 0111111101=> 
 	 	 	 	 <= 00733B
 	 	 	when 0111111110=> 
 	 	 	 	 <= 509G78
 	 	 	when 1000000000=> 
 	 	 	 	 <= E3F6EE
 	 	 	when 1000000001=> 
 	 	 	 	 <= 00733B
 	 	 	when 1000000010=> 
 	 	 	 	 <= 78B688
 	 	 	when 1000000011=> 
 	 	 	 	 <= F47373
 	 	 	when 1000000100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000000101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000000110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000000111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000001000=> 
 	 	 	 	 <= EE6768
 	 	 	when 1000001001=> 
 	 	 	 	 <= 8F4243
 	 	 	when 1000001010=> 
 	 	 	 	 <= DB5G5G
 	 	 	when 1000001011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000001100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000001101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000001110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000001111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000010000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000010001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000010010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000010011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000010100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000010101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000010110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000010111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000011000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000011001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000011010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000011011=> 
 	 	 	 	 <= F16969
 	 	 	when 1000011100=> 
 	 	 	 	 <= CBC5B7
 	 	 	when 1000011101=> 
 	 	 	 	 <= 00733B
 	 	 	when 1000011110=> 
 	 	 	 	 <= 54B17C
 	 	 	when 1000100000=> 
 	 	 	 	 <= F9G3FF
 	 	 	when 1000100001=> 
 	 	 	 	 <= 00733B
 	 	 	when 1000100010=> 
 	 	 	 	 <= 5E9C77
 	 	 	when 1000100011=> 
 	 	 	 	 <= F78080
 	 	 	when 1000100100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000100101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000100110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000100111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000101000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000101001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000101010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000101011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000101100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000101101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000101110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000101111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000110000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000110001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000110010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000110011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000110100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000110101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000110110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000110111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000111000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000111001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000111010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1000111011=> 
 	 	 	 	 <= F16969
 	 	 	when 1000111100=> 
 	 	 	 	 <= B3C6B2
 	 	 	when 1000111101=> 
 	 	 	 	 <= 00733B
 	 	 	when 1000111110=> 
 	 	 	 	 <= 6DBF8E
 	 	 	when 1001000000=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1001000001=> 
 	 	 	 	 <= 087740
 	 	 	when 1001000010=> 
 	 	 	 	 <= 2F8658
 	 	 	when 1001000011=> 
 	 	 	 	 <= FE9798
 	 	 	when 1001000100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001000101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001000110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001000111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001001000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001001001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001001010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001001011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001001100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001001101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001001110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001001111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001010000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001010001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001010010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001010011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001010100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001010101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001010110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001010111=> 
 	 	 	 	 <= F16969
 	 	 	when 1001011000=> 
 	 	 	 	 <= 482222
 	 	 	when 1001011001=> 
 	 	 	 	 <= 622F2F
 	 	 	when 1001011010=> 
 	 	 	 	 <= EG6868
 	 	 	when 1001011011=> 
 	 	 	 	 <= F57676
 	 	 	when 1001011100=> 
 	 	 	 	 <= 75B586
 	 	 	when 1001011101=> 
 	 	 	 	 <= 00733B
 	 	 	when 1001011110=> 
 	 	 	 	 <= 94D4BD
 	 	 	when 1001100001=> 
 	 	 	 	 <= 40966C
 	 	 	when 1001100010=> 
 	 	 	 	 <= 01733B
 	 	 	when 1001100011=> 
 	 	 	 	 <= F7C4C1
 	 	 	when 1001100100=> 
 	 	 	 	 <= F2696B
 	 	 	when 1001100101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001100110=> 
 	 	 	 	 <= F2696B
 	 	 	when 1001100111=> 
 	 	 	 	 <= F1696B
 	 	 	when 1001101000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001101001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001101010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001101011=> 
 	 	 	 	 <= F16969
 	 	 	when 1001101100=> 
 	 	 	 	 <= 9B4848
 	 	 	when 1001101101=> 
 	 	 	 	 <= DD5G60
 	 	 	when 1001101110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001101111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001110000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001110001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001110010=> 
 	 	 	 	 <= 592929
 	 	 	when 1001110011=> 
 	 	 	 	 <= 693131
 	 	 	when 1001110100=> 
 	 	 	 	 <= EF6868
 	 	 	when 1001110101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001110110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1001110111=> 
 	 	 	 	 <= F16969
 	 	 	when 1001111000=> 
 	 	 	 	 <= B04C4C
 	 	 	when 1001111001=> 
 	 	 	 	 <= 562828
 	 	 	when 1001111010=> 
 	 	 	 	 <= EF6868
 	 	 	when 1001111011=> 
 	 	 	 	 <= FE9999
 	 	 	when 1001111100=> 
 	 	 	 	 <= 2F8758
 	 	 	when 1001111101=> 
 	 	 	 	 <= 007339
 	 	 	when 1001111110=> 
 	 	 	 	 <= E0F5EB
 	 	 	when 1010000001=> 
 	 	 	 	 <= 90D2B9
 	 	 	when 1010000010=> 
 	 	 	 	 <= 00733B
 	 	 	when 1010000011=> 
 	 	 	 	 <= 98C29C
 	 	 	when 1010000100=> 
 	 	 	 	 <= F36G70
 	 	 	when 1010000101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010000110=> 
 	 	 	 	 <= 723535
 	 	 	when 1010000111=> 
 	 	 	 	 <= 321717
 	 	 	when 1010001000=> 
 	 	 	 	 <= D65E5E
 	 	 	when 1010001001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010001010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010001011=> 
 	 	 	 	 <= F16969
 	 	 	when 1010001100=> 
 	 	 	 	 <= 572929
 	 	 	when 1010001101=> 
 	 	 	 	 <= 512626
 	 	 	when 1010001110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010001111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010010000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010010001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010010010=> 
 	 	 	 	 <= 9F4B4B
 	 	 	when 1010010011=> 
 	 	 	 	 <= 562828
 	 	 	when 1010010100=> 
 	 	 	 	 <= E36363
 	 	 	when 1010010101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010010110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010010111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010011000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010011001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010011010=> 
 	 	 	 	 <= F16969
 	 	 	when 1010011011=> 
 	 	 	 	 <= E9C8C2
 	 	 	when 1010011100=> 
 	 	 	 	 <= 007239
 	 	 	when 1010011101=> 
 	 	 	 	 <= 157F4B
 	 	 	when 1010011110=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1010100001=> 
 	 	 	 	 <= FDG4G0
 	 	 	when 1010100010=> 
 	 	 	 	 <= 03753D
 	 	 	when 1010100011=> 
 	 	 	 	 <= 258352
 	 	 	when 1010100100=> 
 	 	 	 	 <= FGB4B4
 	 	 	when 1010100101=> 
 	 	 	 	 <= F2696B
 	 	 	when 1010100110=> 
 	 	 	 	 <= E46363
 	 	 	when 1010100111=> 
 	 	 	 	 <= 833E3E
 	 	 	when 1010101000=> 
 	 	 	 	 <= E06161
 	 	 	when 1010101001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010101010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010101011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010101100=> 
 	 	 	 	 <= F16969
 	 	 	when 1010101101=> 
 	 	 	 	 <= F2696B
 	 	 	when 1010101110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010101111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010110000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010110001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010110010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010110011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010110100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010110101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010110110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010110111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010111000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010111001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1010111010=> 
 	 	 	 	 <= F78283
 	 	 	when 1010111011=> 
 	 	 	 	 <= 6CB180
 	 	 	when 1010111100=> 
 	 	 	 	 <= 007239
 	 	 	when 1010111101=> 
 	 	 	 	 <= 77C496
 	 	 	when 1011000010=> 
 	 	 	 	 <= 63B986
 	 	 	when 1011000011=> 
 	 	 	 	 <= 007239
 	 	 	when 1011000100=> 
 	 	 	 	 <= 9EC29E
 	 	 	when 1011000101=> 
 	 	 	 	 <= F47676
 	 	 	when 1011000110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011000111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011001000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011001001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011001010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011001011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011001100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011001101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011001110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011001111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011010000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011010001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011010010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011010011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011010100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011010101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011010110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011010111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011011000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011011001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011011010=> 
 	 	 	 	 <= E7CCC3
 	 	 	when 1011011011=> 
 	 	 	 	 <= 03743D
 	 	 	when 1011011100=> 
 	 	 	 	 <= 06763F
 	 	 	when 1011011101=> 
 	 	 	 	 <= F9G3FF
 	 	 	when 1011100010=> 
 	 	 	 	 <= F8G2FE
 	 	 	when 1011100011=> 
 	 	 	 	 <= 0B7841
 	 	 	when 1011100100=> 
 	 	 	 	 <= 0E7842
 	 	 	when 1011100101=> 
 	 	 	 	 <= EECBC4
 	 	 	when 1011100110=> 
 	 	 	 	 <= F26C6C
 	 	 	when 1011100111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011101000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011101001=> 
 	 	 	 	 <= EE6767
 	 	 	when 1011101010=> 
 	 	 	 	 <= E46363
 	 	 	when 1011101011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011101100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011101101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011101110=> 
 	 	 	 	 <= F16969
 	 	 	when 1011101111=> 
 	 	 	 	 <= 9D4949
 	 	 	when 1011110000=> 
 	 	 	 	 <= E16262
 	 	 	when 1011110001=> 
 	 	 	 	 <= F16969
 	 	 	when 1011110010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011110011=> 
 	 	 	 	 <= F16969
 	 	 	when 1011110100=> 
 	 	 	 	 <= 592929
 	 	 	when 1011110101=> 
 	 	 	 	 <= B14C4C
 	 	 	when 1011110110=> 
 	 	 	 	 <= F1696B
 	 	 	when 1011110111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1011111000=> 
 	 	 	 	 <= F2696B
 	 	 	when 1011111001=> 
 	 	 	 	 <= FFB5B5
 	 	 	when 1011111010=> 
 	 	 	 	 <= 388C5F
 	 	 	when 1011111011=> 
 	 	 	 	 <= 00723B
 	 	 	when 1011111100=> 
 	 	 	 	 <= 7EC79B
 	 	 	when 1011111101=> 
 	 	 	 	 <= GGGFGG
 	 	 	when 1100000011=> 
 	 	 	 	 <= 9DD9C3
 	 	 	when 1100000100=> 
 	 	 	 	 <= 007239
 	 	 	when 1100000101=> 
 	 	 	 	 <= 2E8657
 	 	 	when 1100000110=> 
 	 	 	 	 <= F9C3C0
 	 	 	when 1100000111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1100001000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1100001001=> 
 	 	 	 	 <= 663030
 	 	 	when 1100001010=> 
 	 	 	 	 <= 010000
 	 	 	when 1100001011=> 
 	 	 	 	 <= 8G4343
 	 	 	when 1100001100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1100001101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1100001110=> 
 	 	 	 	 <= EE6868
 	 	 	when 1100001111=> 
 	 	 	 	 <= 431G1G
 	 	 	when 1100010000=> 
 	 	 	 	 <= 5B2B2B
 	 	 	when 1100010001=> 
 	 	 	 	 <= F1696B
 	 	 	when 1100010010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1100010011=> 
 	 	 	 	 <= F16969
 	 	 	when 1100010100=> 
 	 	 	 	 <= 703434
 	 	 	when 1100010101=> 
 	 	 	 	 <= 652G2G
 	 	 	when 1100010110=> 
 	 	 	 	 <= F2696B
 	 	 	when 1100010111=> 
 	 	 	 	 <= F16969
 	 	 	when 1100011000=> 
 	 	 	 	 <= FE9798
 	 	 	when 1100011001=> 
 	 	 	 	 <= 669G7E
 	 	 	when 1100011010=> 
 	 	 	 	 <= 00723B
 	 	 	when 1100011011=> 
 	 	 	 	 <= 298959
 	 	 	when 1100011100=> 
 	 	 	 	 <= GBGDGC
 	 	 	when 1100100011=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1100100100=> 
 	 	 	 	 <= 63B986
 	 	 	when 1100100101=> 
 	 	 	 	 <= 00733B
 	 	 	when 1100100110=> 
 	 	 	 	 <= 33895C
 	 	 	when 1100100111=> 
 	 	 	 	 <= F5C6C3
 	 	 	when 1100101000=> 
 	 	 	 	 <= F36G6G
 	 	 	when 1100101001=> 
 	 	 	 	 <= EC6666
 	 	 	when 1100101010=> 
 	 	 	 	 <= 843F3F
 	 	 	when 1100101011=> 
 	 	 	 	 <= D05B5B
 	 	 	when 1100101100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1100101101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1100101110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1100101111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1100110000=> 
 	 	 	 	 <= F16969
 	 	 	when 1100110001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1100110010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1100110011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1100110100=> 
 	 	 	 	 <= F16969
 	 	 	when 1100110101=> 
 	 	 	 	 <= F2696B
 	 	 	when 1100110110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1100110111=> 
 	 	 	 	 <= FFB3B3
 	 	 	when 1100111000=> 
 	 	 	 	 <= 689G7F
 	 	 	when 1100111001=> 
 	 	 	 	 <= 00733B
 	 	 	when 1100111010=> 
 	 	 	 	 <= 107C46
 	 	 	when 1100111011=> 
 	 	 	 	 <= EFFDF5
 	 	 	when 1101000100=> 
 	 	 	 	 <= GEGFGE
 	 	 	when 1101000101=> 
 	 	 	 	 <= 57B37E
 	 	 	when 1101000110=> 
 	 	 	 	 <= 00733B
 	 	 	when 1101000111=> 
 	 	 	 	 <= 1B7F4C
 	 	 	when 1101001000=> 
 	 	 	 	 <= CGCBBE
 	 	 	when 1101001001=> 
 	 	 	 	 <= FB8G8G
 	 	 	when 1101001010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1101001011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1101001100=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1101001101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1101001110=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1101001111=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1101010000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1101010001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1101010010=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1101010011=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1101010100=> 
 	 	 	 	 <= F2696B
 	 	 	when 1101010101=> 
 	 	 	 	 <= F67E7E
 	 	 	when 1101010110=> 
 	 	 	 	 <= EECBC4
 	 	 	when 1101010111=> 
 	 	 	 	 <= 3E8E62
 	 	 	when 1101011000=> 
 	 	 	 	 <= 007239
 	 	 	when 1101011001=> 
 	 	 	 	 <= 0G7C46
 	 	 	when 1101011010=> 
 	 	 	 	 <= DFF4E9
 	 	 	when 1101100101=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1101100110=> 
 	 	 	 	 <= 7DC799
 	 	 	when 1101100111=> 
 	 	 	 	 <= 00733B
 	 	 	when 1101101000=> 
 	 	 	 	 <= 00723B
 	 	 	when 1101101001=> 
 	 	 	 	 <= 539770
 	 	 	when 1101101010=> 
 	 	 	 	 <= DGCBC1
 	 	 	when 1101101011=> 
 	 	 	 	 <= FF9C9C
 	 	 	when 1101101100=> 
 	 	 	 	 <= F47575
 	 	 	when 1101101101=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1101101110=> 
 	 	 	 	 <= F2696B
 	 	 	when 1101101111=> 
 	 	 	 	 <= F2696B
 	 	 	when 1101110000=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1101110001=> 
 	 	 	 	 <= F26B6B
 	 	 	when 1101110010=> 
 	 	 	 	 <= F36F6F
 	 	 	when 1101110011=> 
 	 	 	 	 <= FC8G8G
 	 	 	when 1101110100=> 
 	 	 	 	 <= F3C6C2
 	 	 	when 1101110101=> 
 	 	 	 	 <= 78B689
 	 	 	when 1101110110=> 
 	 	 	 	 <= 07763F
 	 	 	when 1101110111=> 
 	 	 	 	 <= 00723B
 	 	 	when 1101111000=> 
 	 	 	 	 <= 278858
 	 	 	when 1101111001=> 
 	 	 	 	 <= EEFDF4
 	 	 	when 1110000110=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1110000111=> 
 	 	 	 	 <= D6EGE3
 	 	 	when 1110001000=> 
 	 	 	 	 <= 298959
 	 	 	when 1110001001=> 
 	 	 	 	 <= 00723B
 	 	 	when 1110001010=> 
 	 	 	 	 <= 00723B
 	 	 	when 1110001011=> 
 	 	 	 	 <= 2C8556
 	 	 	when 1110001100=> 
 	 	 	 	 <= 79B789
 	 	 	when 1110001101=> 
 	 	 	 	 <= BGC6B5
 	 	 	when 1110001110=> 
 	 	 	 	 <= DFC5BC
 	 	 	when 1110001111=> 
 	 	 	 	 <= E8C4BE
 	 	 	when 1110010000=> 
 	 	 	 	 <= E3C4BD
 	 	 	when 1110010001=> 
 	 	 	 	 <= CBC6B7
 	 	 	when 1110010010=> 
 	 	 	 	 <= 8DBG95
 	 	 	when 1110010011=> 
 	 	 	 	 <= 439066
 	 	 	when 1110010100=> 
 	 	 	 	 <= 02733C
 	 	 	when 1110010101=> 
 	 	 	 	 <= 00733B
 	 	 	when 1110010110=> 
 	 	 	 	 <= 04753E
 	 	 	when 1110010111=> 
 	 	 	 	 <= 77C496
 	 	 	when 1110011000=> 
 	 	 	 	 <= G9GCGB
 	 	 	when 1110101000=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1110101001=> 
 	 	 	 	 <= BBE0CE
 	 	 	when 1110101010=> 
 	 	 	 	 <= 389266
 	 	 	when 1110101011=> 
 	 	 	 	 <= 00733B
 	 	 	when 1110101100=> 
 	 	 	 	 <= 00733B
 	 	 	when 1110101101=> 
 	 	 	 	 <= 00733B
 	 	 	when 1110101110=> 
 	 	 	 	 <= 007239
 	 	 	when 1110101111=> 
 	 	 	 	 <= 00723B
 	 	 	when 1110110000=> 
 	 	 	 	 <= 00733B
 	 	 	when 1110110001=> 
 	 	 	 	 <= 00733B
 	 	 	when 1110110010=> 
 	 	 	 	 <= 00733B
 	 	 	when 1110110011=> 
 	 	 	 	 <= 00723B
 	 	 	when 1110110100=> 
 	 	 	 	 <= 117D47
 	 	 	when 1110110101=> 
 	 	 	 	 <= 72C192
 	 	 	when 1110110110=> 
 	 	 	 	 <= F6G1FC
 	 	 	when 1110110111=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1111001010=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1111001011=> 
 	 	 	 	 <= FBG3FF
 	 	 	when 1111001100=> 
 	 	 	 	 <= B6DFCB
 	 	 	when 1111001101=> 
 	 	 	 	 <= 74C294
 	 	 	when 1111001110=> 
 	 	 	 	 <= 56B27D
 	 	 	when 1111001111=> 
 	 	 	 	 <= 499C72
 	 	 	when 1111010000=> 
 	 	 	 	 <= 4F9F76
 	 	 	when 1111010001=> 
 	 	 	 	 <= 64B987
 	 	 	when 1111010010=> 
 	 	 	 	 <= 8ED0B7
 	 	 	when 1111010011=> 
 	 	 	 	 <= DBF2E6
 	 	 	when 1111010100=> 
 	 	 	 	 <= GEGFGF 
 	 	 end case; 
     	 end if;  
     end process; 
 address <= row & col; 
 end;
