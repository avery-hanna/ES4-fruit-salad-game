library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ROM is
  port(
	  row : in std_logic_vector(4 downto 0);
	  col : in std_logic_vector(4 downto 0);
	  fruit_color : in std_logic_vector(5 downto 0);
	  clk : in std_logic;
	  color : out std_logic_vector(5 downto 0)
  );
end ROM;

architecture synth of ROM is 
signal address : std_logic_vector(9 downto 0);
begin
	process(clk) is
	begin
		if rising_edge(clk) then
			case address is 

 	 	 	when "0000001100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0000001101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0000001110" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0000001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0000010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0000010001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0000010010" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0000010011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0000101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0000101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0000101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0000101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0000101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0000101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0000110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0000110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0000110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0000110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0000110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0000110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0000110110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0001001000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001001001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001001010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001100101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0001100110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0001100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0001111001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0001111010" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0010000100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0010000101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010000110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010000111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010001000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010001001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010001010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010011010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010011011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0010100011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0010100100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0010111100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0011000011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0011000100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011000101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011000110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011000111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011001000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011001001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011001010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011011100" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0011100011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0011111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100000010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100000011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100000100" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0100000101" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0100000110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100000111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100001000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100001001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100001010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100011010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100011011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100011100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100011101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100100001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0100100010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100100011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100100100" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0100100101" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0100100110" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0100100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100101010" => 
 	 	 	 	 color <= "000110";
 	 	 	when "0100101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0100111110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0101000001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101000010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101000011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101000100" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0101000101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0101000110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0101000111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101001000" => 
 	 	 	 	 color <= "000110";
 	 	 	when "0101001001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0101001010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0101001011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0101001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101011010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101011011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101011100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101011101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101011110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101100001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101100010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101100011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101100100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0101100101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0101100110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0101100111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0101101000" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0101101001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0101101010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0101101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0101111110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110000000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0110000001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110000010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110000011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110000100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0110000101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0110000110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0110000111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0110001000" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0110001001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0110001010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0110001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110011010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110011011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110011100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110011101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110011110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110100000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0110100001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110100010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110100011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0110100100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0110100101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0110100110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0110100111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0110101000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0110101001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0110101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0110111110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111000000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111000001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111000010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0111000011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0111000100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0111000101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0111000110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0111000111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0111001000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0111001001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111001010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111011010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111011011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111011100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111011101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111011110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111100000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111100001" => 
 	 	 	 	 color <= "000110";
 	 	 	when "0111100010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "0111100011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0111100100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0111100101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0111100110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0111100111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0111101000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0111101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "0111111110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000000000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000000001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000000010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000000011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1000000100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1000000101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1000000110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1000000111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1000001000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1000001001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000001010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000011010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000011011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000011100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000011101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000011110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000100000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000100001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000100010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000100011" => 
 	 	 	 	 color <= "000110";
 	 	 	when "1000100100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1000100101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1000100110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1000100111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1000101000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1000101001" => 
 	 	 	 	 color <= "000110";
 	 	 	when "1000101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1000111110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001000000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1001000001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001000010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001000011" => 
 	 	 	 	 color <= "000110";
 	 	 	when "1001000100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1001000101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1001000110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1001000111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1001001000" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1001001001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1001001010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001011010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001011011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001011100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001011101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001011110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001100000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1001100001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001100010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001100011" => 
 	 	 	 	 color <= "000110";
 	 	 	when "1001100100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1001100101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1001100110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1001100111" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1001101000" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1001101001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1001101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1001111110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000011" => 
 	 	 	 	 color <= "000110";
 	 	 	when "1010000100" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010000101" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010000110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010000111" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010001000" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010001001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010001010" => 
 	 	 	 	 color <= "000110";
 	 	 	when "1010001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010011110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100100" => 
 	 	 	 	 color <= "000110";
 	 	 	when "1010100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101000" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010101001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1010101010" => 
 	 	 	 	 color <= "000110";
 	 	 	when "1010101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1010111110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011000010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011000111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "1011001010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011011110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1011100010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1011111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100000010" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1100000011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100000100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100000101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100000110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100000111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100001000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100001001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100001010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100011010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100011011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100011100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100011101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1100100011" => 
 	 	 	 	 color <= "000110";
 	 	 	when "1100100100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1100111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101000011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1101000100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101000101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101000110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101000111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101001000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101001001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101001010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101011010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101011011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101011100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1101100100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1101100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1101111011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1110000101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1110000110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110000111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110001000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110001001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110001010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110011010" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1110100111" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1110101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110101111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1110111000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1111001001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "1111001010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1111001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1111001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1111001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1111001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1111001111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1111010000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1111010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1111010010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1111010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1111010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1111010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "1111010110" => 
 	 	 	 	 color <= "000001"; 
 	 	 end case; 
     	 end if;  
     end process; 
 address <= row & col; 
 end;