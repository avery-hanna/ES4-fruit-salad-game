library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity fruitROM is
  port(
	  row : in std_logic_vector(3 downto 0);
	  col : in std_logic_vector(3 downto 0);
	  fruit_type : in std_logic_vector(2 downto 0);
	  clk : in std_logic;
	  color : out std_logic_vector(5 downto 0)
  );
end fruitROM;

architecture synth of fruitROM is 

signal address: std_logic_vector(10 downto 0);
signal color3: std_logic_vector(2 downto 0);

begin
	process(clk) is
	begin
		if rising_edge(clk) then
			case address is
				--blueberry
				when "00000000101" => 
 	 				color3 <= "00" 
				when "00000000110" => 
					color3 <= "010" 
				when "00000000111" => 
					color3 <= "010" 
				when "00000001000" => 
					color3 <= "010" 
				when "00000001001" => 
					color3 <= "011" 
				when "00000010011" => 
					color3 <= "00" 
				when "00000010100" => 
					color3 <= "010" 
				when "00000010101" => 
					color3 <= "010" 
				when "00000010110" => 
					color3 <= "010" 
				when "00000010111" => 
					color3 <= "010" 
				when "00000011000" => 
					color3 <= "010" 
				when "00000011001" => 
					color3 <= "010" 
				when "00000011010" => 
					color3 <= "010" 
				when "00000011011" => 
					color3 <= "010" 
				when "00000100010" => 
					color3 <= "010" 
				when "00000100011" => 
					color3 <= "010" 
				when "00000100100" => 
					color3 <= "010" 
				when "00000100101" => 
					color3 <= "010" 
				when "00000100110" => 
					color3 <= "010" 
				when "00000100111" => 
					color3 <= "010" 
				when "00000101000" => 
					color3 <= "010" 
				when "00000101001" => 
					color3 <= "010" 
				when "00000101010" => 
					color3 <= "010" 
				when "00000101011" => 
					color3 <= "010" 
				when "00000101100" => 
					color3 <= "010" 
				when "00000110001" => 
					color3 <= "011" 
				when "00000110010" => 
					color3 <= "010" 
				when "00000110011" => 
					color3 <= "010" 
				when "00000110100" => 
					color3 <= "010" 
				when "00000110101" => 
					color3 <= "010" 
				when "00000110110" => 
					color3 <= "010" 
				when "00000110111" => 
					color3 <= "010" 
				when "00000111000" => 
					color3 <= "010" 
				when "00000111001" => 
					color3 <= "010" 
				when "00000111010" => 
					color3 <= "010" 
				when "00000111011" => 
					color3 <= "010" 
				when "00000111100" => 
					color3 <= "010" 
				when "00000111101" => 
					color3 <= "010" 
				when "00000111110" => 
					color3 <= "101" 
				when "00001000001" => 
					color3 <= "010" 
				when "00001000010" => 
					color3 <= "011" 
				when "00001000011" => 
					color3 <= "010" 
				when "00001000100" => 
					color3 <= "010" 
				when "00001000101" => 
					color3 <= "010" 
				when "00001000110" => 
					color3 <= "010" 
				when "00001000111" => 
					color3 <= "010" 
				when "00001001000" => 
					color3 <= "010" 
				when "00001001001" => 
					color3 <= "010" 
				when "00001001010" => 
					color3 <= "010" 
				when "00001001011" => 
					color3 <= "010" 
				when "00001001100" => 
					color3 <= "010" 
				when "00001001101" => 
					color3 <= "010" 
				when "00001001110" => 
					color3 <= "00" 
				when "00001010000" => 
					color3 <= "00" 
				when "00001010001" => 
					color3 <= "010" 
				when "00001010010" => 
					color3 <= "00" 
				when "00001010011" => 
					color3 <= "00" 
				when "00001010100" => 
					color3 <= "011" 
				when "00001010101" => 
					color3 <= "010" 
				when "00001010110" => 
					color3 <= "010" 
				when "00001010111" => 
					color3 <= "010" 
				when "00001011000" => 
					color3 <= "010" 
				when "00001011001" => 
					color3 <= "010" 
				when "00001011010" => 
					color3 <= "010" 
				when "00001011011" => 
					color3 <= "010" 
				when "00001011100" => 
					color3 <= "010" 
				when "00001011101" => 
					color3 <= "010" 
				when "00001011110" => 
					color3 <= "010" 
				when "00001100000" => 
					color3 <= "010" 
				when "00001100001" => 
					color3 <= "100" 
				when "00001100010" => 
					color3 <= "00" 
				when "00001100011" => 
					color3 <= "00" 
				when "00001100100" => 
					color3 <= "011" 
				when "00001100101" => 
					color3 <= "010" 
				when "00001100110" => 
					color3 <= "010" 
				when "00001100111" => 
					color3 <= "010" 
				when "00001101000" => 
					color3 <= "010" 
				when "00001101001" => 
					color3 <= "010" 
				when "00001101010" => 
					color3 <= "010" 
				when "00001101011" => 
					color3 <= "010" 
				when "00001101100" => 
					color3 <= "010" 
				when "00001101101" => 
					color3 <= "010" 
				when "00001101110" => 
					color3 <= "010" 
				when "00001110000" => 
					color3 <= "010" 
				when "00001110001" => 
					color3 <= "00" 
				when "00001110010" => 
					color3 <= "00" 
				when "00001110011" => 
					color3 <= "00" 
				when "00001110100" => 
					color3 <= "010" 
				when "00001110101" => 
					color3 <= "010" 
				when "00001110110" => 
					color3 <= "010" 
				when "00001110111" => 
					color3 <= "010" 
				when "00001111000" => 
					color3 <= "010" 
				when "00001111001" => 
					color3 <= "010" 
				when "00001111010" => 
					color3 <= "010" 
				when "00001111011" => 
					color3 <= "010" 
				when "00001111100" => 
					color3 <= "010" 
				when "00001111101" => 
					color3 <= "010" 
				when "00001111110" => 
					color3 <= "010" 
				when "00010000000" => 
					color3 <= "010" 
				when "00010000001" => 
					color3 <= "010" 
				when "00010000010" => 
					color3 <= "00" 
				when "00010000011" => 
					color3 <= "00" 
				when "00010000100" => 
					color3 <= "100" 
				when "00010000101" => 
					color3 <= "010" 
				when "00010000110" => 
					color3 <= "010" 
				when "00010000111" => 
					color3 <= "010" 
				when "00010001000" => 
					color3 <= "010" 
				when "00010001001" => 
					color3 <= "010" 
				when "00010001010" => 
					color3 <= "010" 
				when "00010001011" => 
					color3 <= "010" 
				when "00010001100" => 
					color3 <= "010" 
				when "00010001101" => 
					color3 <= "010" 
				when "00010001110" => 
					color3 <= "010" 
				when "00010010000" => 
					color3 <= "011" 
				when "00010010001" => 
					color3 <= "010" 
				when "00010010010" => 
					color3 <= "00" 
				when "00010010011" => 
					color3 <= "011" 
				when "00010010100" => 
					color3 <= "011" 
				when "00010010101" => 
					color3 <= "010" 
				when "00010010110" => 
					color3 <= "010" 
				when "00010010111" => 
					color3 <= "010" 
				when "00010011000" => 
					color3 <= "010" 
				when "00010011001" => 
					color3 <= "010" 
				when "00010011010" => 
					color3 <= "010" 
				when "00010011011" => 
					color3 <= "010" 
				when "00010011100" => 
					color3 <= "010" 
				when "00010011101" => 
					color3 <= "010" 
				when "00010011110" => 
					color3 <= "010" 
				when "00010100000" => 
					color3 <= "00" 
				when "00010100001" => 
					color3 <= "010" 
				when "00010100010" => 
					color3 <= "010" 
				when "00010100011" => 
					color3 <= "010" 
				when "00010100100" => 
					color3 <= "011" 
				when "00010100101" => 
					color3 <= "010" 
				when "00010100110" => 
					color3 <= "010" 
				when "00010100111" => 
					color3 <= "010" 
				when "00010101000" => 
					color3 <= "010" 
				when "00010101001" => 
					color3 <= "010" 
				when "00010101010" => 
					color3 <= "010" 
				when "00010101011" => 
					color3 <= "010" 
				when "00010101100" => 
					color3 <= "010" 
				when "00010101101" => 
					color3 <= "010" 
				when "00010101110" => 
					color3 <= "100" 
				when "00010110001" => 
					color3 <= "010" 
				when "00010110010" => 
					color3 <= "010" 
				when "00010110011" => 
					color3 <= "010" 
				when "00010110100" => 
					color3 <= "010" 
				when "00010110101" => 
					color3 <= "010" 
				when "00010110110" => 
					color3 <= "010" 
				when "00010110111" => 
					color3 <= "010" 
				when "00010111000" => 
					color3 <= "010" 
				when "00010111001" => 
					color3 <= "010" 
				when "00010111010" => 
					color3 <= "010" 
				when "00010111011" => 
					color3 <= "010" 
				when "00010111100" => 
					color3 <= "010" 
				when "00010111101" => 
					color3 <= "010" 
				when "00010111110" => 
					color3 <= "101" 
				when "00011000010" => 
					color3 <= "010" 
				when "00011000011" => 
					color3 <= "010" 
				when "00011000100" => 
					color3 <= "010" 
				when "00011000101" => 
					color3 <= "010" 
				when "00011000110" => 
					color3 <= "010" 
				when "00011000111" => 
					color3 <= "010" 
				when "00011001000" => 
					color3 <= "010" 
				when "00011001001" => 
					color3 <= "010" 
				when "00011001010" => 
					color3 <= "010" 
				when "00011001011" => 
					color3 <= "010" 
				when "00011001100" => 
					color3 <= "010" 
				when "00011001101" => 
					color3 <= "00" 
				when "00011010011" => 
					color3 <= "010" 
				when "00011010100" => 
					color3 <= "010" 
				when "00011010101" => 
					color3 <= "010" 
				when "00011010110" => 
					color3 <= "010" 
				when "00011010111" => 
					color3 <= "010" 
				when "00011011000" => 
					color3 <= "010" 
				when "00011011001" => 
					color3 <= "010" 
				when "00011011010" => 
					color3 <= "010" 
				when "00011011011" => 
					color3 <= "010" 
				when "00011011100" => 
					color3 <= "00" 
				when "00011100011" => 
					color3 <= "101" 
				when "00011100100" => 
					color3 <= "00" 
				when "00011100101" => 
					color3 <= "010" 
				when "00011100110" => 
					color3 <= "010" 
				when "00011100111" => 
					color3 <= "010" 
				when "00011101000" => 
					color3 <= "010" 
				when "00011101001" => 
					color3 <= "010" 
				when "00011101010" => 
					color3 <= "100" 
				when "00011101011" => 
					color3 <= "101" 
				--cherry 
				when "00100000101" => 
 	 				color3 <= "001" 
				when "00100000110" => 
					color3 <= "010" 
				when "00100000111" => 
					color3 <= "010" 
				when "00100001000" => 
					color3 <= "010" 
				when "00100001001" => 
					color3 <= "001" 
				when "00100010011" => 
					color3 <= "001" 
				when "00100010100" => 
					color3 <= "010" 
				when "00100010101" => 
					color3 <= "010" 
				when "00100010110" => 
					color3 <= "010" 
				when "00100010111" => 
					color3 <= "010" 
				when "00100011000" => 
					color3 <= "010" 
				when "00100011001" => 
					color3 <= "010" 
				when "00100011010" => 
					color3 <= "010" 
				when "00100011011" => 
					color3 <= "001" 
				when "00100100010" => 
					color3 <= "010" 
				when "00100100011" => 
					color3 <= "010" 
				when "00100100100" => 
					color3 <= "010" 
				when "00100100101" => 
					color3 <= "010" 
				when "00100100110" => 
					color3 <= "010" 
				when "00100100111" => 
					color3 <= "010" 
				when "00100101000" => 
					color3 <= "010" 
				when "00100101001" => 
					color3 <= "010" 
				when "00100101010" => 
					color3 <= "010" 
				when "00100101011" => 
					color3 <= "010" 
				when "00100101100" => 
					color3 <= "010" 
				when "00100110001" => 
					color3 <= "001" 
				when "00100110010" => 
					color3 <= "010" 
				when "00100110011" => 
					color3 <= "010" 
				when "00100110100" => 
					color3 <= "010" 
				when "00100110101" => 
					color3 <= "010" 
				when "00100110110" => 
					color3 <= "010" 
				when "00100110111" => 
					color3 <= "010" 
				when "00100111000" => 
					color3 <= "010" 
				when "00100111001" => 
					color3 <= "010" 
				when "00100111010" => 
					color3 <= "010" 
				when "00100111011" => 
					color3 <= "010" 
				when "00100111100" => 
					color3 <= "010" 
				when "00100111101" => 
					color3 <= "001" 
				when "00101000001" => 
					color3 <= "010" 
				when "00101000001" => 
					color3 <= "010" 
				when "00101000011" => 
					color3 <= "010" 
				when "00101000100" => 
					color3 <= "010" 
				when "00101000101" => 
					color3 <= "010" 
				when "00101000110" => 
					color3 <= "010" 
				when "00101000111" => 
					color3 <= "010" 
				when "00101001000" => 
					color3 <= "010" 
				when "00101001001" => 
					color3 <= "010" 
				when "00101001010" => 
					color3 <= "010" 
				when "00101001011" => 
					color3 <= "010" 
				when "00101001100" => 
					color3 <= "010" 
				when "00101001101" => 
					color3 <= "010" 
				when "00101001110" => 
					color3 <= "101" 
				when "00101010000" => 
					color3 <= "001" 
				when "00101010001" => 
					color3 <= "110" 
				when "00101010010" => 
					color3 <= "111" 
				when "00101010011" => 
					color3 <= "010" 
				when "00101010100" => 
					color3 <= "010" 
				when "00101010101" => 
					color3 <= "010" 
				when "00101010110" => 
					color3 <= "010" 
				when "00101010111" => 
					color3 <= "010" 
				when "00101011000" => 
					color3 <= "010" 
				when "00101011001" => 
					color3 <= "010" 
				when "00101011010" => 
					color3 <= "010" 
				when "00101011011" => 
					color3 <= "010" 
				when "00101011100" => 
					color3 <= "010" 
				when "00101011101" => 
					color3 <= "010" 
				when "00101011110" => 
					color3 <= "001" 
				when "00101100000" => 
					color3 <= "001" 
				when "00101100001" => 
					color3 <= "010" 
				when "00101100010" => 
					color3 <= "110" 
				when "00101100010" => 
					color3 <= "110" 
				when "00101100100" => 
					color3 <= "010" 
				when "00101100101" => 
					color3 <= "010" 
				when "00101100110" => 
					color3 <= "010" 
				when "00101100111" => 
					color3 <= "010" 
				when "00101101000" => 
					color3 <= "010" 
				when "00101101001" => 
					color3 <= "010" 
				when "00101101010" => 
					color3 <= "010" 
				when "00101101011" => 
					color3 <= "010" 
				when "00101101100" => 
					color3 <= "010" 
				when "00101101101" => 
					color3 <= "010" 
				when "00101101110" => 
					color3 <= "010" 
				when "00101110000" => 
					color3 <= "010" 
				when "00101110001" => 
					color3 <= "010" 
				when "00101110010" => 
					color3 <= "011" 
				when "00101110011" => 
					color3 <= "110" 
				when "00101110100" => 
					color3 <= "010" 
				when "00101110101" => 
					color3 <= "010" 
				when "00101110110" => 
					color3 <= "010" 
				when "00101110111" => 
					color3 <= "010" 
				when "00101111000" => 
					color3 <= "010" 
				when "00101111001" => 
					color3 <= "010" 
				when "00101111010" => 
					color3 <= "010" 
				when "00101111011" => 
					color3 <= "010" 
				when "00101111100" => 
					color3 <= "010" 
				when "00101111101" => 
					color3 <= "010" 
				when "00101111110" => 
					color3 <= "010" 
				when "00110000000" => 
					color3 <= "001" 
				when "00110000001" => 
					color3 <= "001" 
				when "00110000010" => 
					color3 <= "011" 
				when "00110000011" => 
					color3 <= "110" 
				when "00110000100" => 
					color3 <= "010" 
				when "00110000101" => 
					color3 <= "010" 
				when "00110000110" => 
					color3 <= "010" 
				when "00110000111" => 
					color3 <= "010" 
				when "00110001000" => 
					color3 <= "010" 
				when "00110001001" => 
					color3 <= "010" 
				when "00110001010" => 
					color3 <= "010" 
				when "00110001011" => 
					color3 <= "010" 
				when "00110001100" => 
					color3 <= "010" 
				when "00110001101" => 
					color3 <= "010" 
				when "00110001110" => 
					color3 <= "010" 
				when "00110010000" => 
					color3 <= "001" 
				when "00110010001" => 
					color3 <= "010" 
				when "00110010010" => 
					color3 <= "010" 
				when "00110010010" => 
					color3 <= "010" 
				when "00110010100" => 
					color3 <= "110" 
				when "00110010101" => 
					color3 <= "111" 
				when "00110010110" => 
					color3 <= "010" 
				when "00110010111" => 
					color3 <= "010" 
				when "00110011000" => 
					color3 <= "010" 
				when "00110011001" => 
					color3 <= "010" 
				when "00110011010" => 
					color3 <= "010" 
				when "00110011011" => 
					color3 <= "010" 
				when "00110011100" => 
					color3 <= "010" 
				when "00110011101" => 
					color3 <= "010" 
				when "00110011110" => 
					color3 <= "010" 
				when "00110100001" => 
					color3 <= "010" 
				when "00110100010" => 
					color3 <= "100" 
				when "00110100011" => 
					color3 <= "010" 
				when "00110100100" => 
					color3 <= "111" 
				when "00110100101" => 
					color3 <= "111" 
				when "00110100101" => 
					color3 <= "111" 
				when "00110100111" => 
					color3 <= "010" 
				when "00110101000" => 
					color3 <= "010" 
				when "00110101001" => 
					color3 <= "010" 
				when "00110101010" => 
					color3 <= "010" 
				when "00110101011" => 
					color3 <= "010" 
				when "00110101100" => 
					color3 <= "010" 
				when "00110101101" => 
					color3 <= "010" 
				when "00110101110" => 
					color3 <= "001" 
				when "00110110001" => 
					color3 <= "010" 
				when "00110110010" => 
					color3 <= "010" 
				when "00110110010" => 
					color3 <= "010" 
				when "00110110100" => 
					color3 <= "111" 
				when "00110110101" => 
					color3 <= "111" 
				when "00110110101" => 
					color3 <= "111" 
				when "00110110111" => 
					color3 <= "010" 
				when "00110111000" => 
					color3 <= "010" 
				when "00110111001" => 
					color3 <= "010" 
				when "00110111010" => 
					color3 <= "010" 
				when "00110111011" => 
					color3 <= "010" 
				when "00110111100" => 
					color3 <= "010" 
				when "00110111101" => 
					color3 <= "010" 
				when "00110111110" => 
					color3 <= "101" 
				when "00111000010" => 
					color3 <= "010" 
				when "00111000011" 
				=> 	 color3 <= "100" 
				when "00111000100" => 
					color3 <= "111" 
				when "00111000100" => 
					color3 <= "111" 
				when "00111000110" => 
					color3 <= "010" 
				when "00111000111" => 
					color3 <= "010" 
				when "00111001000" => 
					color3 <= "010" 
				when "00111001001" => 
					color3 <= "010" 
				when "00111001010" => 
					color3 <= "010" 
				when "00111001011" => 
					color3 <= "010" 
				when "00111001100" => 
					color3 <= "010" 
				when "00111001101" => 
					color3 <= "101" 
				when "00111010011" => 
					color3 <= "010" 
				when "00111010100" => 
					color3 <= "010" 
				when "00111010101" => 
					color3 <= "010" 
				when "00111010110" => 
					color3 <= "010" 
				when "00111010111" => 
					color3 <= "010" 
				when "00111011000" => 
					color3 <= "010" 
				when "00111011001" => 
					color3 <= "010" 
				when "00111011010" => 
					color3 <= "010" 
				when "00111011011" => 
					color3 <= "010" 
				when "00111011100" => 
					color3 <= "101" 
				when "00111100011" => 
					color3 <= "101" 
				when "00111100100" => 
					color3 <= "001" 
				when "00111100101" => 
					color3 <= "010" 
				when "00111100110" => 
					color3 <= "010" 
				when "00111100111" => 
					color3 <= "010" 
				when "00111101000" => 
					color3 <= "010" 
				when "00111101001" => 
					color3 <= "010" 
				when "00111101010" => 
					color3 <= "001" 
				when "00111101011" => 
					color3 <= "101" 
				--watermelon
				when "01000000101" => 
					color3 <= "100" 
				when "01000000110" => 
					color3 <= "110" 
				when "01000000111" => 
					color3 <= "111" 
				when "01000001000" => 
					color3 <= "110" 
				when "01000001001" => 
					color3 <= "111" 
				when "01000010011" => 
					color3 <= "111" 
				when "01000010100" => 
					color3 <= "101" 
				when "01000010101" => 
					color3 <= "011" 
				when "01000010110" => 
					color3 <= "011" 
				when "01000010110" => 
					color3 <= "011" 
				when "01000011000" => 
					color3 <= "011" 
				when "01000011001" => 
					color3 <= "011" 
				when "01000011010" => 
					color3 <= "101" 
				when "01000011011" => 
					color3 <= "111" 
				when "01000100010" => 
					color3 <= "110" 
				when "01000100011" => 
					color3 <= "011" 
				when "01000100011" => 
					color3 <= "011" 
				when "01000100101" => 
					color3 <= "010" 
				when "01000100110" => 
					color3 <= "001" 
				when "01000100111" => 
					color3 <= "001" 
				when "01000101000" => 
					color3 <= "010" 
				when "01000101001" => 
					color3 <= "001" 
				when "01000101001" => 
					color3 <= "001" 
				when "01000101011" => 
					color3 <= "011" 
				when "01000101100" => 
					color3 <= "111" 
				when "01000110001" => 
					color3 <= "111" 
				when "01000110010" => 
					color3 <= "011" 
				when "01000110011" => 
					color3 <= "001" 
				when "01000110100" => 
					color3 <= "010" 
				when "01000110101" => 
					color3 <= "001" 
				when "01000110110" => 
					color3 <= "001" 
				when "01000110111" => 
					color3 <= "001" 
				when "01000111000" => 
					color3 <= "001" 
				when "01000111001" => 
					color3 <= "001" 
				when "01000111010" => 
					color3 <= "010" 
				when "01000111011" => 
					color3 <= "010" 
				when "01000111100" => 
					color3 <= "011" 
				when "01000111101" => 
					color3 <= "110" 
				when "01000111110"=> 
					color3 <= "111" 
				when "01001000001" => 
					color3 <= "101" 
				when "01001000001" => 
					color3 <= "101" 
				when "01001000011" => 
					color3 <= "001" 
				when "01001000100" => 
					color3 <= "010" 
				when "01001000101" => 
					color3 <= "001" 
				when "01001000110" => 
					color3 <= "010" 
				when "01001000111" => 
					color3 <= "010" 
				when "01001001000" => 
					color3 <= "001" 
				when "01001001001" => 
					color3 <= "001" 
				when "01001001010" => 
					color3 <= "010" 
				when "01001001011" => 
					color3 <= "001" 
				when "01001001100" => 
					color3 <= "001" 
				when "01001001101" => 
					color3 <= "101" 
				when "01001001110" => 
					color3 <= "100" 
				when "01001010000" => 
					color3 <= "100" 
				when "01001010001" => 
					color3 <= "011" 
				when "01001010010" => 
					color3 <= "010" 
				when "01001010011" => 
					color3 <= "010" 
				when "01001010100" => 
					color3 <= "010" 
				when "01001010101" => 
					color3 <= "001" 
				when "01001010110" => 
					color3 <= "001" 
				when "01001010111" => 
					color3 <= "001" 
				when "01001011000" => 
					color3 <= "001" 
				when "01001011001" => 
					color3 <= "001" 
				when "01001011010" => 
					color3 <= "001" 
				when "01001011011" => 
					color3 <= "010" 
				when "01001011100" => 
					color3 <= "001" 
				when "01001011101" => 
					color3 <= "011" 
				when "01001011110" => 
					color3 <= "110" 
				when "01001100000" => 
					color3 <= "111" 
				when "01001100001" => 
					color3 <= "011" 
				when "01001100010" => 
					color3 <= "001" 
				when "01001100011" => 
					color3 <= "001" 
				when "01001100100" => 
					color3 <= "001" 
				when "01001100101" => 
					color3 <= "001" 
				when "01001100110" => 
					color3 <= "010" 
				when "01001100111" => 
					color3 <= "001" 
				when "01001101000" => 
					color3 <= "010" 
				when "01001101001" => 
					color3 <= "001" 
				when "01001101010" => 
					color3 <= "001" 
				when "01001101011" => 
					color3 <= "010" 
				when "01001101100" => 
					color3 <= "001" 
				when "01001101100" => 
					color3 <= "001" 
				when "01001101110" => 
					color3 <= "111" 
				when "01001110000" => 
					color3 <= "110" 
				when "01001110000" => 
					color3 <= "110" 
				when "01001110010" => 
					color3 <= "001" 
				when "01001110011" => 
					color3 <= "010" 
				when "01001110100" => 
					color3 <= "001" 
				when "01001110101" => 
					color3 <= "001" 
				when "01001110110" => 
					color3 <= "001" 
				when "01001110111" => 
					color3 <= "001" 
				when "01001111000" => 
					color3 <= "001" 
				when "01001111001" => 
					color3 <= "001" 
				when "01001111010" => 
					color3 <= "010" 
				when "01001111011" => 
					color3 <= "001" 
				when "01001111100" => 
					color3 <= "010" 
				when "01001111100" => 
					color3 <= "010" 
				when "01001111110" => 
					color3 <= "101" 
				when "01010000000" => 
					color3 <= "110" 
				when "01010000001" => 
					color3 <= "011" 
				when "01010000010" => 
					color3 <= "010" 
				when "01010000011" => 
					color3 <= "001" 
				when "01010000100" => 
					color3 <= "001" 
				when "01010000101" => 
					color3 <= "001" 
				when "01010000110" => 
					color3 <= "010" 
				when "01010000111" => 
					color3 <= "001" 
				when "01010001000" => 
					color3 <= "010" 
				when "01010001001" => 
					color3 <= "001" 
				when "01010001010" => 
					color3 <= "001" 
				when "01010001011" => 
					color3 <= "001" 
				when "01010001100" => 
					color3 <= "001" 
				when "01010001100" => 
					color3 <= "001" 
				when "01010001110" => 
					color3 <= "101" 
				when "01010010000" => 
					color3 <= "100" 
				when "01010010001" => 
					color3 <= "011" 
				when "01010010010" => 
					color3 <= "001" 
				when "01010010011" => 
					color3 <= "001" 
				when "01010010100" => 
					color3 <= "010" 
				when "01010010101" => 
					color3 <= "001" 
				when "01010010110" => 
					color3 <= "001" 
				when "01010010111" => 
					color3 <= "001" 
				when "01010011000" => 
					color3 <= "001" 
				when "01010011001" => 
					color3 <= "001" 
				when "01010011010" => 
					color3 <= "001" 
				when "01010011011" => 
					color3 <= "010" 
				when "01010011100" => 
					color3 <= "001" 
				when "01010011101" => 
					color3 <= "011" 
				when "01010011110" => 
					color3 <= "110" 
				when "01010100001" => 
					color3 <= "101" 
				when "01010100001" => 
					color3 <= "101" 
				when "01010100011" => 
					color3 <= "001" 
				when "01010100100" => 
					color3 <= "001" 
				when "01010100101" => 
					color3 <= "001" 
				when "01010100110" => 
					color3 <= "001" 
				when "01010100111" => 
					color3 <= "010" 
				when "01010101000" => 
					color3 <= "010" 
				when "01010101001" => 
					color3 <= "001" 
				when "01010101010" => 
					color3 <= "010" 
				when "01010101011" => 
					color3 <= "001" 
				when "01010101100" => 
					color3 <= "001" 
				when "01010101101" => 
					color3 <= "101" 
				when "01010101110" => 
					color3 <= "100" 
				when "01010110001" => 
					color3 <= "111" 
				when "01010110010" => 
					color3 <= "011" 
				when "01010110011" => 
					color3 <= "001" 
				when "01010110100" => 
					color3 <= "010" 
				when "01010110101" => 
					color3 <= "010" 
				when "01010110110" => 
					color3 <= "001" 
				when "01010110111" => 
					color3 <= "001" 
				when "01010111000" => 
					color3 <= "001" 
				when "01010111001" => 
					color3 <= "001" 
				when "01010111010" => 
					color3 <= "001" 
				when "01010111011" => 
					color3 <= "010" 
				when "01010111100" => 
					color3 <= "011" 
				when "01010111101" => 
					color3 <= "111" 
				when "01010111110"=> 
					color3 <= "111" 
				when "01011000010" => 
					color3 <= "111" 
				when "01011000011" => 
					color3 <= "011" 
				when "01011000011" => 
					color3 <= "011" 
				when "01011000101" => 
					color3 <= "001" 
				when "01011000110" => 
					color3 <= "001" 
				when "01011000111" => 
					color3 <= "010" 
				when "01011001000" => 
					color3 <= "001" 
				when "01011001001" => 
					color3 <= "010" 
				when "01011001010" => 
					color3 <= "001" 
				when "01011001011" => 
					color3 <= "011" 
				when "01011001100" => 
					color3 <= "111" 
				when "01011001101"=> 
					color3 <= "111" 
				when "01011010011" => 
					color3 <= "110" 
				when "01011010100" => 
					color3 <= "101" 
				when "01011010101" => 
					color3 <= "011" 
				when "01011010101" => 
					color3 <= "011" 
				when "01011010101" => 
					color3 <= "011" 
				when "01011010101" => 
					color3 <= "011" 
				when "01011011001" => 
					color3 <= "011" 
				when "01011011010" => 
					color3 <= "101" 
				when "01011011011" => 
					color3 <= "111" 
				when "01011011100"=> 
					color3 <= "111" 
				when "01011100011"=> 
					color3 <= "111" 
				when "01011100100" => 
					color3 <= "100" 
				when "01011100101" => 
					color3 <= "111" 
				when "01011100110" => 
					color3 <= "111" 
				when "01011100111" => 
					color3 <= "101" 
				when "01011101000" => 
					color3 <= "111" 
				when "01011101001" => 
					color3 <= "110" 
				when "01011101010" => 
					color3 <= "100" 
				when "01011101011"=> 
					color3 <= "111" 
				when others
					color3 <= "000"
				end case;
			end if;
	end process;
	address <= fruit_type & row & col

	--blueberry
	color <= "000001" when (fruit_type="000" and color3="001")
	else "010110" when (fruit_type="000" and color3="010")
	else "000101" when (fruit_type="000" and color3="011")
	else "000110" when (fruit_type="000" and color3="100")
	else "010101" when (fruit_type="000" and color3="101")
	--cherry
	else "010000" when (fruit_type="010" and color3="001")
	else "100000" when (fruit_type="010" and color3 = "010")
	else "100100" when (fruit_type="010" and color3 = "011")
	else "110101" when (fruit_type="010" and color3 = "100")
	else "010101" when (fruit_type="010" and color3 = "101")
	else "111010" when (fruit_type="010" and color3 = "110")
	else "111111" when (fruit_type="010" and color3 = "111")
	--watermelon
	else "110001" when (fruit_type="010" and color3="001")
	else "100000" when (fruit_type="010" and color3 = "010")
	else "111001" when (fruit_type="010" and color3 = "011")
	else "000100" when (fruit_type="010" and color3 = "100")
	else "101001" when (fruit_type="010" and color3 = "101")
	else "011000" when (fruit_type="010" and color3 = "110")
	else "011001" when (fruit_type="010" and color3 = "111")
	else "000000"

end;