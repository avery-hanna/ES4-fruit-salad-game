library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ROM is
  port(
	  row : in std_logic_vector(4 downto 0);
	  col : in std_logic_vector(4 downto 0);
	  fruit_color : in std_logic_vector(5 downto 0);
	  clk : in std_logic;
	  color : out std_logic_vector(5 downto 0)
  );
end ROM;

architecture synth of ROM is 
signal address : std_logic_vector(9 downto 0);
begin
	process(clk) is
	begin
		if rising_edge(clk) then
			case address is 

 	 	 	when "0000000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000001001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000100011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0000100100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000100111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0000101011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0001100010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001100111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0001101101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0010000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010001110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0010100000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0010100001" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0010100010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0010100011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010100111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010101000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010101001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010101010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010101011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010101100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010101101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0010101110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0011000000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0011000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011000010" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0011000011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0011000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011001101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011001110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011100000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011100001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011100010" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0011100011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0011100100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011100101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011100110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011100111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011101000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011101001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011101010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011101011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011101100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011101101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0011101110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100000000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100000001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "0100000010" => 
 	 	 	 	 color <= "100100";
 	 	 	when "0100000011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0100000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100001101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100001110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100100000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0100100001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100100010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100100011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0100100100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "0100100101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0100100110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100100111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100101000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100101001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100101010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100101011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100101100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100101101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0100101110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101000010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "0101000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101000100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101000110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101001101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101001110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0101100001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101100010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101100011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101100101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0101100110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0101100111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101101000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101101001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101101010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101101011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101101100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101101101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0101101110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0110000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110000011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "0110000100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "0110000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "0110000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110001101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0110100011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110100100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110100101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110100110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110100111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110101000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110101001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110101010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110101011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0110101100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0111000011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "0111000100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0111000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0111000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0111001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0111001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "0111001010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "0111001011" => 
 	 	 	 	 color <= "000001"; 
 	 	 end case; 
     	 end if;  
     end process; 
 address <= row & col; 
 end;