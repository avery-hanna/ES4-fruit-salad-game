library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity BLUEBERRYROM is
  port(
	  row : in std_logic_vector(4 downto 0);
	  col : in std_logic_vector(4 downto 0);
	  fruit_color : in std_logic_vector(5 downto 0);
	  clk : in std_logic;
	  color : out std_logic_vector(5 downto 0)
  );
end BLUEBERRYROM;

architecture synth of BLUEBERRYROM is 
signal address : std_logic_vector(9 downto 0);
begin
	process(clk) is
	begin
		if rising_edge(clk) then
			case address is 

 	 	 	when 0000001010=> 
 	 	 	 	 <= GEGEGF
 	 	 	when 0000001011=> 
 	 	 	 	 <= E3E6FC
 	 	 	when 0000001100=> 
 	 	 	 	 <= B1B6E5
 	 	 	when 0000001101=> 
 	 	 	 	 <= 7E84D5
 	 	 	when 0000001110=> 
 	 	 	 	 <= 666GCC
 	 	 	when 0000001111=> 
 	 	 	 	 <= 5D65C7
 	 	 	when 0000010000=> 
 	 	 	 	 <= 5E66C7
 	 	 	when 0000010001=> 
 	 	 	 	 <= 6B72CE
 	 	 	when 0000010010=> 
 	 	 	 	 <= 8B91DC
 	 	 	when 0000010011=> 
 	 	 	 	 <= C5C9EF
 	 	 	when 0000010100=> 
 	 	 	 	 <= FDFEG6
 	 	 	when 0000101000=> 
 	 	 	 	 <= G2G2G9
 	 	 	when 0000101001=> 
 	 	 	 	 <= 9DB2E3
 	 	 	when 0000101010=> 
 	 	 	 	 <= 505BC2
 	 	 	when 0000101011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0000101100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0000101101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0000101110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0000101111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0000110000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0000110001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0000110010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0000110011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0000110100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0000110101=> 
 	 	 	 	 <= 6F76CG
 	 	 	when 0000110110=> 
 	 	 	 	 <= D7DCF6
 	 	 	when 0000110111=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0001000110=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0001000111=> 
 	 	 	 	 <= BCBGE9
 	 	 	when 0001001000=> 
 	 	 	 	 <= 4B54BG
 	 	 	when 0001001001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001001010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001001011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001001100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001001101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001001110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001001111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001010000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001010001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001010010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001010011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001010100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001010101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001010110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001010111=> 
 	 	 	 	 <= 6972CD
 	 	 	when 0001011000=> 
 	 	 	 	 <= F0F1G1
 	 	 	when 0001100101=> 
 	 	 	 	 <= G2G3G9
 	 	 	when 0001100110=> 
 	 	 	 	 <= 6G78CG
 	 	 	when 0001100111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001101000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001101001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001101010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001101011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001101100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001101101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001101110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001101111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001110000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001110001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001110010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001110011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001110100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001110101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001110110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001110111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0001111000=> 
 	 	 	 	 <= 4650BE
 	 	 	when 0001111001=> 
 	 	 	 	 <= C2C7EE
 	 	 	when 0010000100=> 
 	 	 	 	 <= FCFDG6
 	 	 	when 0010000101=> 
 	 	 	 	 <= 5B64C6
 	 	 	when 0010000110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010000111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010001000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010001001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010001010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010001011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010001100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010001101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010001110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010001111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010010000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010010001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010010010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010010011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010010100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010010101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010010110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010010111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010011000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010011001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010011010=> 
 	 	 	 	 <= 9CB1E2
 	 	 	when 0010011011=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0010100011=> 
 	 	 	 	 <= G4G4GB
 	 	 	when 0010100100=> 
 	 	 	 	 <= 5D66C7
 	 	 	when 0010100101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010100110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010100111=> 
 	 	 	 	 <= 3E46B6
 	 	 	when 0010101000=> 
 	 	 	 	 <= 2G3097
 	 	 	when 0010101001=> 
 	 	 	 	 <= 3F47B7
 	 	 	when 0010101010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010101011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010101100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010101101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010101110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010101111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010110000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010110001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010110010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010110011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010110100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010110101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010110110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010110111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010111000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010111001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010111010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0010111011=> 
 	 	 	 	 <= B5BBE7
 	 	 	when 0011000010=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0011000011=> 
 	 	 	 	 <= 767FD2
 	 	 	when 0011000100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011000101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011000110=> 
 	 	 	 	 <= 32359B
 	 	 	when 0011000111=> 
 	 	 	 	 <= 120376
 	 	 	when 0011001000=> 
 	 	 	 	 <= 120376
 	 	 	when 0011001001=> 
 	 	 	 	 <= 1D1381
 	 	 	when 0011001010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011001011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011001100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011001101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011001110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011001111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011010000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011010001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011010010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011010011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011010100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011010101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011010110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011010111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011011000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011011001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011011010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011011011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011011100=> 
 	 	 	 	 <= DDDGF8
 	 	 	when 0011100010=> 
 	 	 	 	 <= C7CCEG
 	 	 	when 0011100011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011100100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011100101=> 
 	 	 	 	 <= 33369C
 	 	 	when 0011100110=> 
 	 	 	 	 <= 120376
 	 	 	when 0011100111=> 
 	 	 	 	 <= 120376
 	 	 	when 0011101000=> 
 	 	 	 	 <= 120376
 	 	 	when 0011101001=> 
 	 	 	 	 <= 120376
 	 	 	when 0011101010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011101011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011101100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011101101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011101110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011101111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011110000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011110001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011110010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011110011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011110100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011110101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011110110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011110111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011111000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011111001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011111010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011111011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0011111100=> 
 	 	 	 	 <= 535EC3
 	 	 	when 0011111101=> 
 	 	 	 	 <= G7G8GC
 	 	 	when 0100000001=> 
 	 	 	 	 <= G9GBGD
 	 	 	when 0100000010=> 
 	 	 	 	 <= 505BC1
 	 	 	when 0100000011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100000100=> 
 	 	 	 	 <= 3G49B8
 	 	 	when 0100000101=> 
 	 	 	 	 <= 150779
 	 	 	when 0100000110=> 
 	 	 	 	 <= 120376
 	 	 	when 0100000111=> 
 	 	 	 	 <= 120376
 	 	 	when 0100001000=> 
 	 	 	 	 <= 120376
 	 	 	when 0100001001=> 
 	 	 	 	 <= 110275
 	 	 	when 0100001010=> 
 	 	 	 	 <= 2C2991
 	 	 	when 0100001011=> 
 	 	 	 	 <= 323499
 	 	 	when 0100001100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100001101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100001110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100001111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100010000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100010001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100010010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100010011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100010100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100010101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100010110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100010111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100011000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100011001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100011010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100011011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100011100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100011101=> 
 	 	 	 	 <= 9EB3E4
 	 	 	when 0100100001=> 
 	 	 	 	 <= BGC4EC
 	 	 	when 0100100010=> 
 	 	 	 	 <= 383EB0
 	 	 	when 0100100011=> 
 	 	 	 	 <= 180E7E
 	 	 	when 0100100100=> 
 	 	 	 	 <= 241G8B
 	 	 	when 0100100101=> 
 	 	 	 	 <= 120376
 	 	 	when 0100100110=> 
 	 	 	 	 <= 120376
 	 	 	when 0100100111=> 
 	 	 	 	 <= 130577
 	 	 	when 0100101000=> 
 	 	 	 	 <= 140678
 	 	 	when 0100101001=> 
 	 	 	 	 <= 120376
 	 	 	when 0100101010=> 
 	 	 	 	 <= 120376
 	 	 	when 0100101011=> 
 	 	 	 	 <= 120376
 	 	 	when 0100101100=> 
 	 	 	 	 <= 3C42B3
 	 	 	when 0100101101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100101110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100101111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100110000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100110001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100110010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100110011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100110100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100110101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100110110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100110111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100111000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100111001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100111010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100111011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100111100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0100111101=> 
 	 	 	 	 <= 4C55BG
 	 	 	when 0100111110=> 
 	 	 	 	 <= G8G8GD
 	 	 	when 0101000000=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0101000001=> 
 	 	 	 	 <= 5G68C8
 	 	 	when 0101000010=> 
 	 	 	 	 <= 160B7C
 	 	 	when 0101000011=> 
 	 	 	 	 <= 120376
 	 	 	when 0101000100=> 
 	 	 	 	 <= 120376
 	 	 	when 0101000101=> 
 	 	 	 	 <= 120376
 	 	 	when 0101000110=> 
 	 	 	 	 <= 120376
 	 	 	when 0101000111=> 
 	 	 	 	 <= 313298
 	 	 	when 0101001000=> 
 	 	 	 	 <= 150779
 	 	 	when 0101001001=> 
 	 	 	 	 <= 120376
 	 	 	when 0101001010=> 
 	 	 	 	 <= 120376
 	 	 	when 0101001011=> 
 	 	 	 	 <= 120376
 	 	 	when 0101001100=> 
 	 	 	 	 <= 2B2890
 	 	 	when 0101001101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101001110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101001111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101010000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101010001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101010010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101010011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101010100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101010101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101010110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101010111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101011000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101011001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101011010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101011011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101011100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101011101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101011110=> 
 	 	 	 	 <= C8CDF0
 	 	 	when 0101100000=> 
 	 	 	 	 <= F9FBG5
 	 	 	when 0101100001=> 
 	 	 	 	 <= 35399E
 	 	 	when 0101100010=> 
 	 	 	 	 <= 120376
 	 	 	when 0101100011=> 
 	 	 	 	 <= 120376
 	 	 	when 0101100100=> 
 	 	 	 	 <= 120376
 	 	 	when 0101100101=> 
 	 	 	 	 <= 120376
 	 	 	when 0101100110=> 
 	 	 	 	 <= 1B107G
 	 	 	when 0101100111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101101000=> 
 	 	 	 	 <= 16097B
 	 	 	when 0101101001=> 
 	 	 	 	 <= 120376
 	 	 	when 0101101010=> 
 	 	 	 	 <= 120376
 	 	 	when 0101101011=> 
 	 	 	 	 <= 120376
 	 	 	when 0101101100=> 
 	 	 	 	 <= 303297
 	 	 	when 0101101101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101101110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101101111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101110000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101110001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101110010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101110011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101110100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101110101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101110110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101110111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101111000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101111001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101111010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101111011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101111100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101111101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0101111110=> 
 	 	 	 	 <= 7B81D4
 	 	 	when 0110000000=> 
 	 	 	 	 <= C9CEF0
 	 	 	when 0110000001=> 
 	 	 	 	 <= 303197
 	 	 	when 0110000010=> 
 	 	 	 	 <= 120376
 	 	 	when 0110000011=> 
 	 	 	 	 <= 120376
 	 	 	when 0110000100=> 
 	 	 	 	 <= 150779
 	 	 	when 0110000101=> 
 	 	 	 	 <= 190F7F
 	 	 	when 0110000110=> 
 	 	 	 	 <= 373D9G
 	 	 	when 0110000111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110001000=> 
 	 	 	 	 <= 35389D
 	 	 	when 0110001001=> 
 	 	 	 	 <= 1B107G
 	 	 	when 0110001010=> 
 	 	 	 	 <= 120376
 	 	 	when 0110001011=> 
 	 	 	 	 <= 120376
 	 	 	when 0110001100=> 
 	 	 	 	 <= 4049B9
 	 	 	when 0110001101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110001110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110001111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110010000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110010001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110010010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110010011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110010100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110010101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110010110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110010111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110011000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110011001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110011010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110011011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110011100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110011101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110011110=> 
 	 	 	 	 <= 4D56C0
 	 	 	when 0110100000=> 
 	 	 	 	 <= 969DE0
 	 	 	when 0110100001=> 
 	 	 	 	 <= 313399
 	 	 	when 0110100010=> 
 	 	 	 	 <= 120376
 	 	 	when 0110100011=> 
 	 	 	 	 <= 120376
 	 	 	when 0110100100=> 
 	 	 	 	 <= 363B9E
 	 	 	when 0110100101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110100110=> 
 	 	 	 	 <= 414CBB
 	 	 	when 0110100111=> 
 	 	 	 	 <= 414DBB
 	 	 	when 0110101000=> 
 	 	 	 	 <= 3E45B5
 	 	 	when 0110101001=> 
 	 	 	 	 <= 140678
 	 	 	when 0110101010=> 
 	 	 	 	 <= 120376
 	 	 	when 0110101011=> 
 	 	 	 	 <= 130578
 	 	 	when 0110101100=> 
 	 	 	 	 <= 3C42B3
 	 	 	when 0110101101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110101110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110101111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110110000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110110001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110110010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110110011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110110100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110110101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110110110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110110111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110111000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110111001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110111010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110111011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110111100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110111101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0110111110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111000000=> 
 	 	 	 	 <= 8289D7
 	 	 	when 0111000001=> 
 	 	 	 	 <= 383EB0
 	 	 	when 0111000010=> 
 	 	 	 	 <= 120376
 	 	 	when 0111000011=> 
 	 	 	 	 <= 120376
 	 	 	when 0111000100=> 
 	 	 	 	 <= 180D7D
 	 	 	when 0111000101=> 
 	 	 	 	 <= 3F46B6
 	 	 	when 0111000110=> 
 	 	 	 	 <= 27238E
 	 	 	when 0111000111=> 
 	 	 	 	 <= 2D2C93
 	 	 	when 0111001000=> 
 	 	 	 	 <= 26228D
 	 	 	when 0111001001=> 
 	 	 	 	 <= 120376
 	 	 	when 0111001010=> 
 	 	 	 	 <= 120376
 	 	 	when 0111001011=> 
 	 	 	 	 <= 120376
 	 	 	when 0111001100=> 
 	 	 	 	 <= 1C1080
 	 	 	when 0111001101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111001110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111001111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111010000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111010001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111010010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111010011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111010100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111010101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111010110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111010111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111011000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111011001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111011010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111011011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111011100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111011101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111011110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111100000=> 
 	 	 	 	 <= 7B82D4
 	 	 	when 0111100001=> 
 	 	 	 	 <= 424DBC
 	 	 	when 0111100010=> 
 	 	 	 	 <= 140678
 	 	 	when 0111100011=> 
 	 	 	 	 <= 120376
 	 	 	when 0111100100=> 
 	 	 	 	 <= 120376
 	 	 	when 0111100101=> 
 	 	 	 	 <= 34389D
 	 	 	when 0111100110=> 
 	 	 	 	 <= 1G1885
 	 	 	when 0111100111=> 
 	 	 	 	 <= 26218D
 	 	 	when 0111101000=> 
 	 	 	 	 <= 34369C
 	 	 	when 0111101001=> 
 	 	 	 	 <= 110375
 	 	 	when 0111101010=> 
 	 	 	 	 <= 120376
 	 	 	when 0111101011=> 
 	 	 	 	 <= 120376
 	 	 	when 0111101100=> 
 	 	 	 	 <= 120376
 	 	 	when 0111101101=> 
 	 	 	 	 <= 3D43B4
 	 	 	when 0111101110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111101111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111110000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111110001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111110010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111110011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111110100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111110101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111110110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111110111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111111000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111111001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111111010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111111011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111111100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111111101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 0111111110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000000000=> 
 	 	 	 	 <= 7G87D6
 	 	 	when 1000000001=> 
 	 	 	 	 <= 25218C
 	 	 	when 1000000010=> 
 	 	 	 	 <= 120376
 	 	 	when 1000000011=> 
 	 	 	 	 <= 120376
 	 	 	when 1000000100=> 
 	 	 	 	 <= 160B7C
 	 	 	when 1000000101=> 
 	 	 	 	 <= 414CB9
 	 	 	when 1000000110=> 
 	 	 	 	 <= 241F89
 	 	 	when 1000000111=> 
 	 	 	 	 <= 1G1885
 	 	 	when 1000001000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000001001=> 
 	 	 	 	 <= 211B87
 	 	 	when 1000001010=> 
 	 	 	 	 <= 120376
 	 	 	when 1000001011=> 
 	 	 	 	 <= 120376
 	 	 	when 1000001100=> 
 	 	 	 	 <= 120376
 	 	 	when 1000001101=> 
 	 	 	 	 <= 2G2G96
 	 	 	when 1000001110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000001111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000010000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000010001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000010010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000010011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000010100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000010101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000010110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000010111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000011000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000011001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000011010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000011011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000011100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000011101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000011110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000100000=> 
 	 	 	 	 <= 9298DF
 	 	 	when 1000100001=> 
 	 	 	 	 <= 231F89
 	 	 	when 1000100010=> 
 	 	 	 	 <= 120376
 	 	 	when 1000100011=> 
 	 	 	 	 <= 120376
 	 	 	when 1000100100=> 
 	 	 	 	 <= 120376
 	 	 	when 1000100101=> 
 	 	 	 	 <= 1D1381
 	 	 	when 1000100110=> 
 	 	 	 	 <= 383EB0
 	 	 	when 1000100111=> 
 	 	 	 	 <= 383EB0
 	 	 	when 1000101000=> 
 	 	 	 	 <= 424EBC
 	 	 	when 1000101001=> 
 	 	 	 	 <= 190F7F
 	 	 	when 1000101010=> 
 	 	 	 	 <= 120376
 	 	 	when 1000101011=> 
 	 	 	 	 <= 120376
 	 	 	when 1000101100=> 
 	 	 	 	 <= 120376
 	 	 	when 1000101101=> 
 	 	 	 	 <= 2F2F95
 	 	 	when 1000101110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000101111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000110000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000110001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000110010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000110011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000110100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000110101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000110110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000110111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000111000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000111001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000111010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000111011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000111100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000111101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1000111110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001000000=> 
 	 	 	 	 <= BGC4ED
 	 	 	when 1001000001=> 
 	 	 	 	 <= 414DBB
 	 	 	when 1001000010=> 
 	 	 	 	 <= 2C2991
 	 	 	when 1001000011=> 
 	 	 	 	 <= 120376
 	 	 	when 1001000100=> 
 	 	 	 	 <= 120376
 	 	 	when 1001000101=> 
 	 	 	 	 <= 120376
 	 	 	when 1001000110=> 
 	 	 	 	 <= 3D44B5
 	 	 	when 1001000111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001001000=> 
 	 	 	 	 <= 3G49B8
 	 	 	when 1001001001=> 
 	 	 	 	 <= 120376
 	 	 	when 1001001010=> 
 	 	 	 	 <= 120376
 	 	 	when 1001001011=> 
 	 	 	 	 <= 120376
 	 	 	when 1001001100=> 
 	 	 	 	 <= 170B7C
 	 	 	when 1001001101=> 
 	 	 	 	 <= 3G49B8
 	 	 	when 1001001110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001001111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001010000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001010001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001010010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001010011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001010100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001010101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001010110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001010111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001011000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001011001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001011010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001011011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001011100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001011101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001011110=> 
 	 	 	 	 <= 4650BE
 	 	 	when 1001100000=> 
 	 	 	 	 <= EDEFFG
 	 	 	when 1001100001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001100010=> 
 	 	 	 	 <= 34389D
 	 	 	when 1001100011=> 
 	 	 	 	 <= 120376
 	 	 	when 1001100100=> 
 	 	 	 	 <= 120376
 	 	 	when 1001100101=> 
 	 	 	 	 <= 120376
 	 	 	when 1001100110=> 
 	 	 	 	 <= 33369B
 	 	 	when 1001100111=> 
 	 	 	 	 <= 424EBC
 	 	 	when 1001101000=> 
 	 	 	 	 <= 3C42B3
 	 	 	when 1001101001=> 
 	 	 	 	 <= 190E7E
 	 	 	when 1001101010=> 
 	 	 	 	 <= 120376
 	 	 	when 1001101011=> 
 	 	 	 	 <= 110275
 	 	 	when 1001101100=> 
 	 	 	 	 <= 3C42B3
 	 	 	when 1001101101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001101110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001101111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001110000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001110001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001110010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001110011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001110100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001110101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001110110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001110111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001111000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001111001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001111010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001111011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001111100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001111101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1001111110=> 
 	 	 	 	 <= 6D74CF
 	 	 	when 1010000000=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1010000001=> 
 	 	 	 	 <= 515CC2
 	 	 	when 1010000010=> 
 	 	 	 	 <= 424EBC
 	 	 	when 1010000011=> 
 	 	 	 	 <= 150879
 	 	 	when 1010000100=> 
 	 	 	 	 <= 120376
 	 	 	when 1010000101=> 
 	 	 	 	 <= 120376
 	 	 	when 1010000110=> 
 	 	 	 	 <= 35399E
 	 	 	when 1010000111=> 
 	 	 	 	 <= 28258F
 	 	 	when 1010001000=> 
 	 	 	 	 <= 120376
 	 	 	when 1010001001=> 
 	 	 	 	 <= 120376
 	 	 	when 1010001010=> 
 	 	 	 	 <= 120376
 	 	 	when 1010001011=> 
 	 	 	 	 <= 120376
 	 	 	when 1010001100=> 
 	 	 	 	 <= 2G3096
 	 	 	when 1010001101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010001110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010001111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010010000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010010001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010010010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010010011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010010100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010010101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010010110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010010111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010011000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010011001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010011010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010011011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010011100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010011101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010011110=> 
 	 	 	 	 <= B7BDE8
 	 	 	when 1010100001=> 
 	 	 	 	 <= 989FE1
 	 	 	when 1010100010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010100011=> 
 	 	 	 	 <= 190F7F
 	 	 	when 1010100100=> 
 	 	 	 	 <= 120376
 	 	 	when 1010100101=> 
 	 	 	 	 <= 120376
 	 	 	when 1010100110=> 
 	 	 	 	 <= 2E2E94
 	 	 	when 1010100111=> 
 	 	 	 	 <= 180D7D
 	 	 	when 1010101000=> 
 	 	 	 	 <= 120376
 	 	 	when 1010101001=> 
 	 	 	 	 <= 120376
 	 	 	when 1010101010=> 
 	 	 	 	 <= 120376
 	 	 	when 1010101011=> 
 	 	 	 	 <= 120376
 	 	 	when 1010101100=> 
 	 	 	 	 <= 29268G
 	 	 	when 1010101101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010101110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010101111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010110000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010110001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010110010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010110011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010110100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010110101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010110110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010110111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010111000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010111001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010111010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010111011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010111100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1010111101=> 
 	 	 	 	 <= 444GBD
 	 	 	when 1010111110=> 
 	 	 	 	 <= FFFGG7
 	 	 	when 1011000001=> 
 	 	 	 	 <= FEFFG7
 	 	 	when 1011000010=> 
 	 	 	 	 <= 4550BE
 	 	 	when 1011000011=> 
 	 	 	 	 <= 25208C
 	 	 	when 1011000100=> 
 	 	 	 	 <= 120376
 	 	 	when 1011000101=> 
 	 	 	 	 <= 120376
 	 	 	when 1011000110=> 
 	 	 	 	 <= 120376
 	 	 	when 1011000111=> 
 	 	 	 	 <= 120376
 	 	 	when 1011001000=> 
 	 	 	 	 <= 120376
 	 	 	when 1011001001=> 
 	 	 	 	 <= 120376
 	 	 	when 1011001010=> 
 	 	 	 	 <= 120376
 	 	 	when 1011001011=> 
 	 	 	 	 <= 120376
 	 	 	when 1011001100=> 
 	 	 	 	 <= 2F2F95
 	 	 	when 1011001101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011001110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011001111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011010000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011010001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011010010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011010011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011010100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011010101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011010110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011010111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011011000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011011001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011011010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011011011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011011100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011011101=> 
 	 	 	 	 <= 868ED9
 	 	 	when 1011100010=> 
 	 	 	 	 <= 989FE1
 	 	 	when 1011100011=> 
 	 	 	 	 <= 3940B2
 	 	 	when 1011100100=> 
 	 	 	 	 <= 120376
 	 	 	when 1011100101=> 
 	 	 	 	 <= 120376
 	 	 	when 1011100110=> 
 	 	 	 	 <= 120376
 	 	 	when 1011100111=> 
 	 	 	 	 <= 120376
 	 	 	when 1011101000=> 
 	 	 	 	 <= 120376
 	 	 	when 1011101001=> 
 	 	 	 	 <= 120376
 	 	 	when 1011101010=> 
 	 	 	 	 <= 120376
 	 	 	when 1011101011=> 
 	 	 	 	 <= 110275
 	 	 	when 1011101100=> 
 	 	 	 	 <= 3D43B4
 	 	 	when 1011101101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011101110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011101111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011110000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011110001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011110010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011110011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011110100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011110101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011110110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011110111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011111000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011111001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011111010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011111011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1011111100=> 
 	 	 	 	 <= 4751BE
 	 	 	when 1011111101=> 
 	 	 	 	 <= F9FBG5
 	 	 	when 1100000010=> 
 	 	 	 	 <= G9G9GD
 	 	 	when 1100000011=> 
 	 	 	 	 <= 5C64C6
 	 	 	when 1100000100=> 
 	 	 	 	 <= 1G1784
 	 	 	when 1100000101=> 
 	 	 	 	 <= 120376
 	 	 	when 1100000110=> 
 	 	 	 	 <= 120376
 	 	 	when 1100000111=> 
 	 	 	 	 <= 1G1784
 	 	 	when 1100001000=> 
 	 	 	 	 <= 120376
 	 	 	when 1100001001=> 
 	 	 	 	 <= 120376
 	 	 	when 1100001010=> 
 	 	 	 	 <= 120376
 	 	 	when 1100001011=> 
 	 	 	 	 <= 1B107G
 	 	 	when 1100001100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100001101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100001110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100001111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100010000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100010001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100010010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100010011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100010100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100010101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100010110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100010111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100011000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100011001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100011010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100011011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100011100=> 
 	 	 	 	 <= BBBGE9
 	 	 	when 1100100011=> 
 	 	 	 	 <= EGF1G1
 	 	 	when 1100100100=> 
 	 	 	 	 <= 4953BF
 	 	 	when 1100100101=> 
 	 	 	 	 <= 33369B
 	 	 	when 1100100110=> 
 	 	 	 	 <= 33369C
 	 	 	when 1100100111=> 
 	 	 	 	 <= 424EBC
 	 	 	when 1100101000=> 
 	 	 	 	 <= 32359B
 	 	 	when 1100101001=> 
 	 	 	 	 <= 1G1784
 	 	 	when 1100101010=> 
 	 	 	 	 <= 221D88
 	 	 	when 1100101011=> 
 	 	 	 	 <= 3C42B3
 	 	 	when 1100101100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100101101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100101110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100101111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100110000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100110001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100110010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100110011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100110100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100110101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100110110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100110111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100111000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100111001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100111010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1100111011=> 
 	 	 	 	 <= 7D84D5
 	 	 	when 1100111100=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1101000100=> 
 	 	 	 	 <= DGE2FB
 	 	 	when 1101000101=> 
 	 	 	 	 <= 4752BF
 	 	 	when 1101000110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101000111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101001000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101001001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101001010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101001011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101001100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101001101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101001110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101001111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101010000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101010001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101010010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101010011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101010100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101010101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101010110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101010111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101011000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101011001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101011010=> 
 	 	 	 	 <= 7078D0
 	 	 	when 1101011011=> 
 	 	 	 	 <= GBGBGD
 	 	 	when 1101100101=> 
 	 	 	 	 <= E7E9FE
 	 	 	when 1101100110=> 
 	 	 	 	 <= 515CC2
 	 	 	when 1101100111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101101000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101101001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101101010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101101011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101101100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101101101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101101110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101101111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101110000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101110001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101110010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101110011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101110100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101110101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101110110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101110111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101111000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1101111001=> 
 	 	 	 	 <= 8188D7
 	 	 	when 1101111010=> 
 	 	 	 	 <= GBGCGE
 	 	 	when 1110000110=> 
 	 	 	 	 <= FGG0G8
 	 	 	when 1110000111=> 
 	 	 	 	 <= 7981D4
 	 	 	when 1110001000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110001001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110001010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110001011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110001100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110001101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110001110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110001111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110010000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110010001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110010010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110010011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110010100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110010101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110010110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110010111=> 
 	 	 	 	 <= 4B55BG
 	 	 	when 1110011000=> 
 	 	 	 	 <= C3C7EE
 	 	 	when 1110101000=> 
 	 	 	 	 <= DEE0F9
 	 	 	when 1110101001=> 
 	 	 	 	 <= 6D75CF
 	 	 	when 1110101010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110101011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110101100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110101101=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110101110=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110101111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110110000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110110001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110110010=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110110011=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110110100=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1110110101=> 
 	 	 	 	 <= 4953BF
 	 	 	when 1110110110=> 
 	 	 	 	 <= 939BDG
 	 	 	when 1110110111=> 
 	 	 	 	 <= G0G1G8
 	 	 	when 1111001010=> 
 	 	 	 	 <= F2F3G2
 	 	 	when 1111001011=> 
 	 	 	 	 <= B1B6E5
 	 	 	when 1111001100=> 
 	 	 	 	 <= 6F77CG
 	 	 	when 1111001101=> 
 	 	 	 	 <= 4B55BG
 	 	 	when 1111001110=> 
 	 	 	 	 <= 424FBD
 	 	 	when 1111001111=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1111010000=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1111010001=> 
 	 	 	 	 <= 434FBD
 	 	 	when 1111010010=> 
 	 	 	 	 <= 5963C5
 	 	 	when 1111010011=> 
 	 	 	 	 <= 838CD8
 	 	 	when 1111010100=> 
 	 	 	 	 <= CDD0F1
 	 	 	when 1111010101=> 
 	 	 	 	 <= G8G8GC 
 	 	 end case; 
     	 end if;  
     end process; 
 address <= row & col; 
 end;
