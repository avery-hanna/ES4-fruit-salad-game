library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity blueberryCherryROM is
  port(
	  fruit_type : in std_logic;
	  row : in std_logic_vector(3 downto 0);
	  col : in std_logic_vector(3 downto 0);
	  clk : in std_logic;
	  color : out std_logic_vector(5 downto 0)
  );
end blueberryCherryROM;

architecture synth of blueberryCherryROM is 
signal address : std_logic_vector(8 downto 0);
begin
	process(clk) is
	begin
		if rising_edge(clk) then
			case address is 

 	 	 	when "000000101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "000000110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000000111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000001000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000001001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "000010011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "000010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000011010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000011011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000100010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000100011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000100100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000110001" => 
 	 	 	 	 color <= "000101";
 	 	 	when "000110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "000111110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "001000001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001000010" => 
 	 	 	 	 color <= "000101";
 	 	 	when "001000011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001000100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001000101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001000110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001000111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001001000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001001001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001001010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001001110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "001010000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "001010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001010010" => 
 	 	 	 	 color <= "000001";
 	 	 	when "001010011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "001010100" => 
 	 	 	 	 color <= "000101";
 	 	 	when "001010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001011010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001011011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001011100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001011101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001011110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001100000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001100001" => 
 	 	 	 	 color <= "000110";
 	 	 	when "001100010" => 
 	 	 	 	 color <= "000001";
 	 	 	when "001100011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "001100100" => 
 	 	 	 	 color <= "000101";
 	 	 	when "001100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001101110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001110000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001110001" => 
 	 	 	 	 color <= "000001";
 	 	 	when "001110010" => 
 	 	 	 	 color <= "000001";
 	 	 	when "001110011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "001110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "001111110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010000000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010000001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010000010" => 
 	 	 	 	 color <= "000001";
 	 	 	when "010000011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "010000100" => 
 	 	 	 	 color <= "000110";
 	 	 	when "010000101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010000110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010000111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010001000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010001001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010001010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010001101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010001110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010010000" => 
 	 	 	 	 color <= "000101";
 	 	 	when "010010001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010010010" => 
 	 	 	 	 color <= "000001";
 	 	 	when "010010011" => 
 	 	 	 	 color <= "000101";
 	 	 	when "010010100" => 
 	 	 	 	 color <= "000101";
 	 	 	when "010010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010011010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010011011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010011100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010011101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010011110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010100000" => 
 	 	 	 	 color <= "000001";
 	 	 	when "010100001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010100010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010100011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010100100" => 
 	 	 	 	 color <= "000101";
 	 	 	when "010100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010101010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010101011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010101100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010101101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010101110" => 
 	 	 	 	 color <= "000110";
 	 	 	when "010110001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010110010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010110011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010110100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010110101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010110110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010110111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010111000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010111001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010111010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010111011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010111100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010111101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "010111110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "011000010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011000011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011000100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011000101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011000110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011000111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011001000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011001001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011001010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011001011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011001100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011001101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "011010011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011010100" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011010101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011010110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011010111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011011000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011011001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011011010" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011011011" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011011100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "011100011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "011100100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "011100101" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011100110" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011100111" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011101000" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011101001" => 
 	 	 	 	 color <= "010110";
 	 	 	when "011101010" => 
 	 	 	 	 color <= "000110";
 	 	 	when "011101011" => 
 	 	 	 	 color <= "000001"; 
			 	 	 	when "100000101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "100000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100001001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "100010011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "100010100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100010101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100010110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100010111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100011000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100011001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100011010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100011011" => 
 	 	 	 	 color <= "010000";
 	 	 	when "100100010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100100011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100100100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100100101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100100110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100100111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100101000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100101001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100101010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100101011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100101100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100110001" => 
 	 	 	 	 color <= "010000";
 	 	 	when "100110010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100110011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100110100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100110101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100110110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100110111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100111000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100111001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100111010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "100111101" => 
 	 	 	 	 color <= "010000";
 	 	 	when "101000001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101000010" => 
 	 	 	 	 color <= "110101";
 	 	 	when "101000011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101001101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101001110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "101010000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "101010001" => 
 	 	 	 	 color <= "111010";
 	 	 	when "101010010" => 
 	 	 	 	 color <= "111111";
 	 	 	when "101010011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101010100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101010101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101010110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101010111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101011000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101011001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101011010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101011011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101011100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101011101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101011110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "101100000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "101100001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101100010" => 
 	 	 	 	 color <= "111010";
 	 	 	when "101100011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "101100100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101100101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101100110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101100111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101101000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101101001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101101010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101101011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101101100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101101101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101101110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101110000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101110001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101110010" => 
 	 	 	 	 color <= "100100";
 	 	 	when "101110011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "101110100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101110101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101110110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101110111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101111000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101111001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101111010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "101111110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110000000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "110000001" => 
 	 	 	 	 color <= "011000";
 	 	 	when "110000010" => 
 	 	 	 	 color <= "100100";
 	 	 	when "110000011" => 
 	 	 	 	 color <= "111010";
 	 	 	when "110000100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110000101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110001101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110001110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110010000" => 
 	 	 	 	 color <= "010000";
 	 	 	when "110010001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110010010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110010011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "110010100" => 
 	 	 	 	 color <= "111010";
 	 	 	when "110010101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "110010110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110010111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110011000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110011001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110011010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110011011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110011100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110011101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110011110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110100001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110100010" => 
 	 	 	 	 color <= "100101";
 	 	 	when "110100011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110100100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "110100101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "110100110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "110100111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110101000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110101001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110101010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110101011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110101100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110101101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110101110" => 
 	 	 	 	 color <= "010000";
 	 	 	when "110110001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110110010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110110011" => 
 	 	 	 	 color <= "110101";
 	 	 	when "110110100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "110110101" => 
 	 	 	 	 color <= "111111";
 	 	 	when "110110110" => 
 	 	 	 	 color <= "110101";
 	 	 	when "110110111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110111000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110111001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110111010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110111011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110111100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110111101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "110111110" => 
 	 	 	 	 color <= "000001";
 	 	 	when "111000010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111000011" => 
 	 	 	 	 color <= "111001";
 	 	 	when "111000100" => 
 	 	 	 	 color <= "111111";
 	 	 	when "111000101" => 
 	 	 	 	 color <= "110101";
 	 	 	when "111000110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111000111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111001000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111001001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111001010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111001011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111001100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111001101" => 
 	 	 	 	 color <= "000001";
 	 	 	when "111010011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111010100" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111010101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111010110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111010111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111011000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111011001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111011010" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111011011" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111011100" => 
 	 	 	 	 color <= "000001";
 	 	 	when "111100011" => 
 	 	 	 	 color <= "000001";
 	 	 	when "111100100" => 
 	 	 	 	 color <= "010000";
 	 	 	when "111100101" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111100110" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111100111" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111101000" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111101001" => 
 	 	 	 	 color <= "100000";
 	 	 	when "111101010" => 
 	 	 	 	 color <= "010000";
 	 	 	when "111101011" => 
 	 	 	 	 color <= "000001";
			when others =>
				color <= "000000";
 	 	 end case;
     	 end if;  
     end process; 
 address <= fruit_type & col & row; 
 end;