library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ROM is
  port(
	  row : in std_logic_vector(4 downto 0);
	  col : in std_logic_vector(4 downto 0);
	  fruit_color : in std_logic_vector(5 downto 0);
	  clk : in std_logic;
	  color : out std_logic_vector(5 downto 0)
  );
end ROM;

architecture synth of ROM is 
signal address : std_logic_vector(9 downto 0);
begin
	process(clk) is
	begin
		if rising_edge(clk) then
			case address is 

 	 	 	when 0000001100=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000001101=> 
 	 	 	 	 <= GFGDG8
 	 	 	when 0000001110=> 
 	 	 	 	 <= GFG2EF
 	 	 	when 0000001111=> 
 	 	 	 	 <= GEFEE0
 	 	 	when 0000010000=> 
 	 	 	 	 <= GFFFE5
 	 	 	when 0000010001=> 
 	 	 	 	 <= GFG7FD
 	 	 	when 0000010010=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000101001=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000101010=> 
 	 	 	 	 <= GEF6CG
 	 	 	when 0000101011=> 
 	 	 	 	 <= GCD364
 	 	 	when 0000101100=> 
 	 	 	 	 <= G9B81G
 	 	 	when 0000101101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0000101110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0000101111=> 
 	 	 	 	 <= G99D00
 	 	 	when 0000110000=> 
 	 	 	 	 <= G99D00
 	 	 	when 0000110001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0000110010=> 
 	 	 	 	 <= G9B009
 	 	 	when 0000110011=> 
 	 	 	 	 <= GBC643
 	 	 	when 0000110100=> 
 	 	 	 	 <= GDE594
 	 	 	when 0000110101=> 
 	 	 	 	 <= GFG8FF
 	 	 	when 0001000111=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0001001000=> 
 	 	 	 	 <= GDEEB9
 	 	 	when 0001001001=> 
 	 	 	 	 <= G9BB23
 	 	 	when 0001001010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0001001011=> 
 	 	 	 	 <= G99F02
 	 	 	when 0001001100=> 
 	 	 	 	 <= GBC02E
 	 	 	when 0001001101=> 
 	 	 	 	 <= GCD257
 	 	 	when 0001001110=> 
 	 	 	 	 <= GDDF70
 	 	 	when 0001001111=> 
 	 	 	 	 <= GDE27B
 	 	 	when 0001010000=> 
 	 	 	 	 <= GDE075
 	 	 	when 0001010001=> 
 	 	 	 	 <= GDD761
 	 	 	when 0001010010=> 
 	 	 	 	 <= GBC73E
 	 	 	when 0001010011=> 
 	 	 	 	 <= G9B20D
 	 	 	when 0001010100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0001010101=> 
 	 	 	 	 <= G99F05
 	 	 	when 0001010110=> 
 	 	 	 	 <= GCD467
 	 	 	when 0001010111=> 
 	 	 	 	 <= GFG7FC
 	 	 	when 0001100101=> 
 	 	 	 	 <= GGGFGF
 	 	 	when 0001100110=> 
 	 	 	 	 <= GFG6F8
 	 	 	when 0001100111=> 
 	 	 	 	 <= GBC53G
 	 	 	when 0001101000=> 
 	 	 	 	 <= G99D00
 	 	 	when 0001101001=> 
 	 	 	 	 <= G9B717
 	 	 	when 0001101010=> 
 	 	 	 	 <= GDDF73
 	 	 	when 0001101011=> 
 	 	 	 	 <= GFFEC8
 	 	 	when 0001101100=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0001101101=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0001101110=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 0001101111=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0001110000=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0001110001=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0001110010=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0001110011=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0001110100=> 
 	 	 	 	 <= GEEC8G
 	 	 	when 0001110101=> 
 	 	 	 	 <= GBC435
 	 	 	when 0001110110=> 
 	 	 	 	 <= G99D00
 	 	 	when 0001110111=> 
 	 	 	 	 <= G9B10D
 	 	 	when 0001111000=> 
 	 	 	 	 <= GDECB3
 	 	 	when 0001111001=> 
 	 	 	 	 <= GFGGGG
 	 	 	when 0010000101=> 
 	 	 	 	 <= GEFCDD
 	 	 	when 0010000110=> 
 	 	 	 	 <= G9B414
 	 	 	when 0010000111=> 
 	 	 	 	 <= G99F03
 	 	 	when 0010001000=> 
 	 	 	 	 <= GDDB68
 	 	 	when 0010001001=> 
 	 	 	 	 <= GFG0CF
 	 	 	when 0010001010=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 0010001011=> 
 	 	 	 	 <= GFF6BB
 	 	 	when 0010001100=> 
 	 	 	 	 <= GDD967
 	 	 	when 0010001101=> 
 	 	 	 	 <= GBC437
 	 	 	when 0010001110=> 
 	 	 	 	 <= G9B819
 	 	 	when 0010001111=> 
 	 	 	 	 <= G9B513
 	 	 	when 0010010000=> 
 	 	 	 	 <= GBBG2B
 	 	 	when 0010010001=> 
 	 	 	 	 <= GDE27C
 	 	 	when 0010010010=> 
 	 	 	 	 <= GFFFCC
 	 	 	when 0010010011=> 
 	 	 	 	 <= GEF2B0
 	 	 	when 0010010100=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0010010101=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 0010010110=> 
 	 	 	 	 <= GEEE93
 	 	 	when 0010010111=> 
 	 	 	 	 <= G9B718
 	 	 	when 0010011000=> 
 	 	 	 	 <= G99D00
 	 	 	when 0010011001=> 
 	 	 	 	 <= GCD66C
 	 	 	when 0010011010=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0010100100=> 
 	 	 	 	 <= GEFBDC
 	 	 	when 0010100101=> 
 	 	 	 	 <= G9B009
 	 	 	when 0010100110=> 
 	 	 	 	 <= G9B411
 	 	 	when 0010100111=> 
 	 	 	 	 <= GEF09C
 	 	 	when 0010101000=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0010101001=> 
 	 	 	 	 <= GFFFCB
 	 	 	when 0010101010=> 
 	 	 	 	 <= GBC73D
 	 	 	when 0010101011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0010101100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0010101101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0010101110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0010101111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0010110000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0010110001=> 
 	 	 	 	 <= GCCF4D
 	 	 	when 0010110010=> 
 	 	 	 	 <= GCD65G
 	 	 	when 0010110011=> 
 	 	 	 	 <= G99D00
 	 	 	when 0010110100=> 
 	 	 	 	 <= G9B81B
 	 	 	when 0010110101=> 
 	 	 	 	 <= GEE582
 	 	 	when 0010110110=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0010110111=> 
 	 	 	 	 <= GFFEC9
 	 	 	when 0010111000=> 
 	 	 	 	 <= GBC538
 	 	 	when 0010111001=> 
 	 	 	 	 <= G89D00
 	 	 	when 0010111010=> 
 	 	 	 	 <= GCD260
 	 	 	when 0010111011=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0011000011=> 
 	 	 	 	 <= GFG5F5
 	 	 	when 0011000100=> 
 	 	 	 	 <= G9B311
 	 	 	when 0011000101=> 
 	 	 	 	 <= G9B411
 	 	 	when 0011000110=> 
 	 	 	 	 <= GFF6B9
 	 	 	when 0011000111=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0011001000=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0011001001=> 
 	 	 	 	 <= GEEC90
 	 	 	when 0011001010=> 
 	 	 	 	 <= G99D00
 	 	 	when 0011001011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011001100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011001101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011001110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011001111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011010000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011010001=> 
 	 	 	 	 <= GDE178
 	 	 	when 0011010010=> 
 	 	 	 	 <= GBC230
 	 	 	when 0011010011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011010100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011010101=> 
 	 	 	 	 <= G99D00
 	 	 	when 0011010110=> 
 	 	 	 	 <= GBC63C
 	 	 	when 0011010111=> 
 	 	 	 	 <= GFFEC8
 	 	 	when 0011011000=> 
 	 	 	 	 <= GFG0CG
 	 	 	when 0011011001=> 
 	 	 	 	 <= GBC73E
 	 	 	when 0011011010=> 
 	 	 	 	 <= G99D00
 	 	 	when 0011011011=> 
 	 	 	 	 <= GDE086
 	 	 	when 0011011100=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0011100010=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0011100011=> 
 	 	 	 	 <= GBC33C
 	 	 	when 0011100100=> 
 	 	 	 	 <= G99F04
 	 	 	when 0011100101=> 
 	 	 	 	 <= GEF19F
 	 	 	when 0011100110=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 0011100111=> 
 	 	 	 	 <= GDDD6F
 	 	 	when 0011101000=> 
 	 	 	 	 <= GBC230
 	 	 	when 0011101001=> 
 	 	 	 	 <= GEF19F
 	 	 	when 0011101010=> 
 	 	 	 	 <= GBC333
 	 	 	when 0011101011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011101100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011101101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011101110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011101111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011110000=> 
 	 	 	 	 <= G99D00
 	 	 	when 0011110001=> 
 	 	 	 	 <= GFF4B4
 	 	 	when 0011110010=> 
 	 	 	 	 <= G9B008
 	 	 	when 0011110011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011110100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011110101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0011110110=> 
 	 	 	 	 <= G89D00
 	 	 	when 0011110111=> 
 	 	 	 	 <= GBBD23
 	 	 	when 0011111000=> 
 	 	 	 	 <= GFFFCB
 	 	 	when 0011111001=> 
 	 	 	 	 <= GFFGCD
 	 	 	when 0011111010=> 
 	 	 	 	 <= GBBD24
 	 	 	when 0011111011=> 
 	 	 	 	 <= G99E01
 	 	 	when 0011111100=> 
 	 	 	 	 <= GEFBDB
 	 	 	when 0100000010=> 
 	 	 	 	 <= GDEDB4
 	 	 	when 0100000011=> 
 	 	 	 	 <= G99D00
 	 	 	when 0100000100=> 
 	 	 	 	 <= GDDC6B
 	 	 	when 0100000101=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 0100000110=> 
 	 	 	 	 <= GDDE6G
 	 	 	when 0100000111=> 
 	 	 	 	 <= G99D00
 	 	 	when 0100001000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100001001=> 
 	 	 	 	 <= G9B615
 	 	 	when 0100001010=> 
 	 	 	 	 <= GFF6B9
 	 	 	when 0100001011=> 
 	 	 	 	 <= G9B30F
 	 	 	when 0100001100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100001101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100001110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100001111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100010000=> 
 	 	 	 	 <= G99G06
 	 	 	when 0100010001=> 
 	 	 	 	 <= GFF4B5
 	 	 	when 0100010010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100010011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100010100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100010101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100010110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100010111=> 
 	 	 	 	 <= G99D00
 	 	 	when 0100011000=> 
 	 	 	 	 <= GEED91
 	 	 	when 0100011001=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0100011010=> 
 	 	 	 	 <= GFF6B8
 	 	 	when 0100011011=> 
 	 	 	 	 <= G99F04
 	 	 	when 0100011100=> 
 	 	 	 	 <= GBBF2D
 	 	 	when 0100011101=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0100100001=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0100100010=> 
 	 	 	 	 <= G9B81G
 	 	 	when 0100100011=> 
 	 	 	 	 <= G9B719
 	 	 	when 0100100100=> 
 	 	 	 	 <= GFG0CG
 	 	 	when 0100100101=> 
 	 	 	 	 <= GFF4B5
 	 	 	when 0100100110=> 
 	 	 	 	 <= G99F03
 	 	 	when 0100100111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100101000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100101001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100101010=> 
 	 	 	 	 <= GCC83G
 	 	 	when 0100101011=> 
 	 	 	 	 <= GEEB8F
 	 	 	when 0100101100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100101101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100101110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100101111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100110000=> 
 	 	 	 	 <= GBC12F
 	 	 	when 0100110001=> 
 	 	 	 	 <= GDE17B
 	 	 	when 0100110010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100110011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100110100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100110101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0100110110=> 
 	 	 	 	 <= G99F03
 	 	 	when 0100110111=> 
 	 	 	 	 <= GDDC6C
 	 	 	when 0100111000=> 
 	 	 	 	 <= GFF8BE
 	 	 	when 0100111001=> 
 	 	 	 	 <= GFFDC5
 	 	 	when 0100111010=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0100111011=> 
 	 	 	 	 <= GCD45B
 	 	 	when 0100111100=> 
 	 	 	 	 <= G99D00
 	 	 	when 0100111101=> 
 	 	 	 	 <= GEF0BG
 	 	 	when 0101000001=> 
 	 	 	 	 <= GEF4C9
 	 	 	when 0101000010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101000011=> 
 	 	 	 	 <= GDE075
 	 	 	when 0101000100=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0101000101=> 
 	 	 	 	 <= GBC538
 	 	 	when 0101000110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101000111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101001000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101001001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101001010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101001011=> 
 	 	 	 	 <= GDE077
 	 	 	when 0101001100=> 
 	 	 	 	 <= GCD357
 	 	 	when 0101001101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101001110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101001111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101010000=> 
 	 	 	 	 <= GCD45C
 	 	 	when 0101010001=> 
 	 	 	 	 <= GCCF4E
 	 	 	when 0101010010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101010011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101010100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101010101=> 
 	 	 	 	 <= GBBC20
 	 	 	when 0101010110=> 
 	 	 	 	 <= GFF2B0
 	 	 	when 0101010111=> 
 	 	 	 	 <= GDD660
 	 	 	when 0101011000=> 
 	 	 	 	 <= G99E02
 	 	 	when 0101011001=> 
 	 	 	 	 <= G99G06
 	 	 	when 0101011010=> 
 	 	 	 	 <= GFFBC3
 	 	 	when 0101011011=> 
 	 	 	 	 <= GFFCC4
 	 	 	when 0101011100=> 
 	 	 	 	 <= G99F03
 	 	 	when 0101011101=> 
 	 	 	 	 <= GBC43E
 	 	 	when 0101011110=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0101100001=> 
 	 	 	 	 <= GCD15F
 	 	 	when 0101100010=> 
 	 	 	 	 <= G99F03
 	 	 	when 0101100011=> 
 	 	 	 	 <= GFFEC9
 	 	 	when 0101100100=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0101100101=> 
 	 	 	 	 <= G9B411
 	 	 	when 0101100110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101100111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101101000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101101001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101101010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101101011=> 
 	 	 	 	 <= G99G05
 	 	 	when 0101101100=> 
 	 	 	 	 <= GFF3B2
 	 	 	when 0101101101=> 
 	 	 	 	 <= GBBD25
 	 	 	when 0101101110=> 
 	 	 	 	 <= G89D00
 	 	 	when 0101101111=> 
 	 	 	 	 <= G89D00
 	 	 	when 0101110000=> 
 	 	 	 	 <= GEE787
 	 	 	when 0101110001=> 
 	 	 	 	 <= GBBC22
 	 	 	when 0101110010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101110011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101110100=> 
 	 	 	 	 <= GCD358
 	 	 	when 0101110101=> 
 	 	 	 	 <= GFF4B4
 	 	 	when 0101110110=> 
 	 	 	 	 <= GBBE26
 	 	 	when 0101110111=> 
 	 	 	 	 <= G99D00
 	 	 	when 0101111000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101111001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101111010=> 
 	 	 	 	 <= GDD762
 	 	 	when 0101111011=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0101111100=> 
 	 	 	 	 <= GBC73D
 	 	 	when 0101111101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0101111110=> 
 	 	 	 	 <= GFG8FE
 	 	 	when 0110000000=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0110000001=> 
 	 	 	 	 <= G9B618
 	 	 	when 0110000010=> 
 	 	 	 	 <= GBC230
 	 	 	when 0110000011=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0110000100=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0110000101=> 
 	 	 	 	 <= GDE47G
 	 	 	when 0110000110=> 
 	 	 	 	 <= GBBE25
 	 	 	when 0110000111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110001000=> 
 	 	 	 	 <= G89D00
 	 	 	when 0110001001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110001010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110001011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110001100=> 
 	 	 	 	 <= GBBC21
 	 	 	when 0110001101=> 
 	 	 	 	 <= GFF4B5
 	 	 	when 0110001110=> 
 	 	 	 	 <= G9B007
 	 	 	when 0110001111=> 
 	 	 	 	 <= G99D00
 	 	 	when 0110010000=> 
 	 	 	 	 <= GFF8BF
 	 	 	when 0110010001=> 
 	 	 	 	 <= G99E01
 	 	 	when 0110010010=> 
 	 	 	 	 <= G9B615
 	 	 	when 0110010011=> 
 	 	 	 	 <= GEEE94
 	 	 	when 0110010100=> 
 	 	 	 	 <= GDDF72
 	 	 	when 0110010101=> 
 	 	 	 	 <= G99G05
 	 	 	when 0110010110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110010111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110011000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110011001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110011010=> 
 	 	 	 	 <= G9B91E
 	 	 	when 0110011011=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0110011100=> 
 	 	 	 	 <= GDE077
 	 	 	when 0110011101=> 
 	 	 	 	 <= G99D00
 	 	 	when 0110011110=> 
 	 	 	 	 <= GDEFBC
 	 	 	when 0110100000=> 
 	 	 	 	 <= GFGBG3
 	 	 	when 0110100001=> 
 	 	 	 	 <= G99D00
 	 	 	when 0110100010=> 
 	 	 	 	 <= GCD45B
 	 	 	when 0110100011=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0110100100=> 
 	 	 	 	 <= GFF9BG
 	 	 	when 0110100101=> 
 	 	 	 	 <= GDE077
 	 	 	when 0110100110=> 
 	 	 	 	 <= GEEB8F
 	 	 	when 0110100111=> 
 	 	 	 	 <= GFF9BG
 	 	 	when 0110101000=> 
 	 	 	 	 <= GEEE94
 	 	 	when 0110101001=> 
 	 	 	 	 <= GDDB68
 	 	 	when 0110101010=> 
 	 	 	 	 <= GBC73D
 	 	 	when 0110101011=> 
 	 	 	 	 <= G9B411
 	 	 	when 0110101100=> 
 	 	 	 	 <= G99D00
 	 	 	when 0110101101=> 
 	 	 	 	 <= GCD359
 	 	 	when 0110101110=> 
 	 	 	 	 <= GEE889
 	 	 	when 0110101111=> 
 	 	 	 	 <= GCCC46
 	 	 	when 0110110000=> 
 	 	 	 	 <= GEF29G
 	 	 	when 0110110001=> 
 	 	 	 	 <= GCCD48
 	 	 	when 0110110010=> 
 	 	 	 	 <= GFF6B9
 	 	 	when 0110110011=> 
 	 	 	 	 <= GBC435
 	 	 	when 0110110100=> 
 	 	 	 	 <= G99D00
 	 	 	when 0110110101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110110110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110110111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110111000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110111001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0110111010=> 
 	 	 	 	 <= G99D00
 	 	 	when 0110111011=> 
 	 	 	 	 <= GFFEC8
 	 	 	when 0110111100=> 
 	 	 	 	 <= GEF3B1
 	 	 	when 0110111101=> 
 	 	 	 	 <= G99D00
 	 	 	when 0110111110=> 
 	 	 	 	 <= GCDC78
 	 	 	when 0111000000=> 
 	 	 	 	 <= GFFFE4
 	 	 	when 0111000001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111000010=> 
 	 	 	 	 <= GDDG75
 	 	 	when 0111000011=> 
 	 	 	 	 <= GGG0D1
 	 	 	when 0111000100=> 
 	 	 	 	 <= GBBG2B
 	 	 	when 0111000101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111000110=> 
 	 	 	 	 <= G99D00
 	 	 	when 0111000111=> 
 	 	 	 	 <= G99D00
 	 	 	when 0111001000=> 
 	 	 	 	 <= G9B514
 	 	 	when 0111001001=> 
 	 	 	 	 <= GCC840
 	 	 	when 0111001010=> 
 	 	 	 	 <= GDDC6D
 	 	 	when 0111001011=> 
 	 	 	 	 <= GEEG98
 	 	 	when 0111001100=> 
 	 	 	 	 <= GFF8BE
 	 	 	when 0111001101=> 
 	 	 	 	 <= GFF6B9
 	 	 	when 0111001110=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0111001111=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0111010000=> 
 	 	 	 	 <= GGG0D1
 	 	 	when 0111010001=> 
 	 	 	 	 <= GEE889
 	 	 	when 0111010010=> 
 	 	 	 	 <= G9B20D
 	 	 	when 0111010011=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111010100=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111010101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111010110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111010111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111011000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111011001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111011010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111011011=> 
 	 	 	 	 <= GEF09D
 	 	 	when 0111011100=> 
 	 	 	 	 <= GFFFCC
 	 	 	when 0111011101=> 
 	 	 	 	 <= G99D00
 	 	 	when 0111011110=> 
 	 	 	 	 <= GCCG58
 	 	 	when 0111100000=> 
 	 	 	 	 <= GEF9D7
 	 	 	when 0111100001=> 
 	 	 	 	 <= G89D00
 	 	 	when 0111100010=> 
 	 	 	 	 <= GDE47G
 	 	 	when 0111100011=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0111100100=> 
 	 	 	 	 <= G9B10B
 	 	 	when 0111100101=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111100110=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111100111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111101000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111101001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111101010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111101011=> 
 	 	 	 	 <= G99D00
 	 	 	when 0111101100=> 
 	 	 	 	 <= G99G06
 	 	 	when 0111101101=> 
 	 	 	 	 <= GDDC6B
 	 	 	when 0111101110=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 0111101111=> 
 	 	 	 	 <= GFG1D0
 	 	 	when 0111110000=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 0111110001=> 
 	 	 	 	 <= GFF6B9
 	 	 	when 0111110010=> 
 	 	 	 	 <= GDE077
 	 	 	when 0111110011=> 
 	 	 	 	 <= GCCE4C
 	 	 	when 0111110100=> 
 	 	 	 	 <= GBBB1G
 	 	 	when 0111110101=> 
 	 	 	 	 <= G99E01
 	 	 	when 0111110110=> 
 	 	 	 	 <= G99D00
 	 	 	when 0111110111=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111111000=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111111001=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111111010=> 
 	 	 	 	 <= G99E00
 	 	 	when 0111111011=> 
 	 	 	 	 <= GEEF97
 	 	 	when 0111111100=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 0111111101=> 
 	 	 	 	 <= G99D00
 	 	 	when 0111111110=> 
 	 	 	 	 <= GBCB4E
 	 	 	when 1000000000=> 
 	 	 	 	 <= GEFCDD
 	 	 	when 1000000001=> 
 	 	 	 	 <= G99D00
 	 	 	when 1000000010=> 
 	 	 	 	 <= GDE27B
 	 	 	when 1000000011=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1000000100=> 
 	 	 	 	 <= G9B30F
 	 	 	when 1000000101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000000110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000000111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000001000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000001001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000001010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000001011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000001100=> 
 	 	 	 	 <= G9B109
 	 	 	when 1000001101=> 
 	 	 	 	 <= GEEF96
 	 	 	when 1000001110=> 
 	 	 	 	 <= GFFEC8
 	 	 	when 1000001111=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1000010000=> 
 	 	 	 	 <= GFFEC8
 	 	 	when 1000010001=> 
 	 	 	 	 <= GBBD25
 	 	 	when 1000010010=> 
 	 	 	 	 <= GBC231
 	 	 	when 1000010011=> 
 	 	 	 	 <= GCD55E
 	 	 	when 1000010100=> 
 	 	 	 	 <= GEE889
 	 	 	when 1000010101=> 
 	 	 	 	 <= GFF9BF
 	 	 	when 1000010110=> 
 	 	 	 	 <= GEEE94
 	 	 	when 1000010111=> 
 	 	 	 	 <= GDDB68
 	 	 	when 1000011000=> 
 	 	 	 	 <= GBC73D
 	 	 	when 1000011001=> 
 	 	 	 	 <= G9B411
 	 	 	when 1000011010=> 
 	 	 	 	 <= G99F02
 	 	 	when 1000011011=> 
 	 	 	 	 <= GFFFCC
 	 	 	when 1000011100=> 
 	 	 	 	 <= GFG0CG
 	 	 	when 1000011101=> 
 	 	 	 	 <= G99D00
 	 	 	when 1000011110=> 
 	 	 	 	 <= GBCC50
 	 	 	when 1000100000=> 
 	 	 	 	 <= GFG3F0
 	 	 	when 1000100001=> 
 	 	 	 	 <= G99D00
 	 	 	when 1000100010=> 
 	 	 	 	 <= GDD967
 	 	 	when 1000100011=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1000100100=> 
 	 	 	 	 <= GBBE25
 	 	 	when 1000100101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000100110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000100111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000101000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000101001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000101010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000101011=> 
 	 	 	 	 <= GBBE26
 	 	 	when 1000101100=> 
 	 	 	 	 <= GFF4B4
 	 	 	when 1000101101=> 
 	 	 	 	 <= GCD359
 	 	 	when 1000101110=> 
 	 	 	 	 <= G9B10C
 	 	 	when 1000101111=> 
 	 	 	 	 <= GFFGCF
 	 	 	when 1000110000=> 
 	 	 	 	 <= GFF5B6
 	 	 	when 1000110001=> 
 	 	 	 	 <= GDDC6B
 	 	 	when 1000110010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000110011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000110100=> 
 	 	 	 	 <= G99D00
 	 	 	when 1000110101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1000110110=> 
 	 	 	 	 <= G9B514
 	 	 	when 1000110111=> 
 	 	 	 	 <= GCC840
 	 	 	when 1000111000=> 
 	 	 	 	 <= GDDC6D
 	 	 	when 1000111001=> 
 	 	 	 	 <= GEEG98
 	 	 	when 1000111010=> 
 	 	 	 	 <= GFFEC8
 	 	 	when 1000111011=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1000111100=> 
 	 	 	 	 <= GFF8BE
 	 	 	when 1000111101=> 
 	 	 	 	 <= G99D00
 	 	 	when 1000111110=> 
 	 	 	 	 <= GCD465
 	 	 	when 1001000000=> 
 	 	 	 	 <= GFGFGE
 	 	 	when 1001000001=> 
 	 	 	 	 <= G99F03
 	 	 	when 1001000010=> 
 	 	 	 	 <= GCCB43
 	 	 	when 1001000011=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1001000100=> 
 	 	 	 	 <= GCCG4F
 	 	 	when 1001000101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001000110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001000111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001001000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001001001=> 
 	 	 	 	 <= G99E01
 	 	 	when 1001001010=> 
 	 	 	 	 <= GDD760
 	 	 	when 1001001011=> 
 	 	 	 	 <= GEF2B0
 	 	 	when 1001001100=> 
 	 	 	 	 <= GBBC20
 	 	 	when 1001001101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001001110=> 
 	 	 	 	 <= GBBB20
 	 	 	when 1001001111=> 
 	 	 	 	 <= GEE889
 	 	 	when 1001010000=> 
 	 	 	 	 <= G99E01
 	 	 	when 1001010001=> 
 	 	 	 	 <= GEEG98
 	 	 	when 1001010010=> 
 	 	 	 	 <= GBC333
 	 	 	when 1001010011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001010100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001010101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001010110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001010111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001011000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001011001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001011010=> 
 	 	 	 	 <= GCCG4F
 	 	 	when 1001011011=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1001011100=> 
 	 	 	 	 <= GEE889
 	 	 	when 1001011101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001011110=> 
 	 	 	 	 <= GDE38F
 	 	 	when 1001100001=> 
 	 	 	 	 <= GBC136
 	 	 	when 1001100010=> 
 	 	 	 	 <= G9B411
 	 	 	when 1001100011=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1001100100=> 
 	 	 	 	 <= GEE98C
 	 	 	when 1001100101=> 
 	 	 	 	 <= G99D00
 	 	 	when 1001100110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001100111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001101000=> 
 	 	 	 	 <= G9B819
 	 	 	when 1001101001=> 
 	 	 	 	 <= GEF09B
 	 	 	when 1001101010=> 
 	 	 	 	 <= GDDC6C
 	 	 	when 1001101011=> 
 	 	 	 	 <= G99F03
 	 	 	when 1001101100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001101101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001101110=> 
 	 	 	 	 <= GCCF4D
 	 	 	when 1001101111=> 
 	 	 	 	 <= GCD55D
 	 	 	when 1001110000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001110001=> 
 	 	 	 	 <= G9B615
 	 	 	when 1001110010=> 
 	 	 	 	 <= GFF6B9
 	 	 	when 1001110011=> 
 	 	 	 	 <= G9B30F
 	 	 	when 1001110100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001110101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001110110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001110111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001111000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001111001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1001111010=> 
 	 	 	 	 <= GCCD49
 	 	 	when 1001111011=> 
 	 	 	 	 <= GGG0D1
 	 	 	when 1001111100=> 
 	 	 	 	 <= GCD155
 	 	 	when 1001111101=> 
 	 	 	 	 <= G99D00
 	 	 	when 1001111110=> 
 	 	 	 	 <= GEFBDB
 	 	 	when 1010000001=> 
 	 	 	 	 <= GDE085
 	 	 	when 1010000010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010000011=> 
 	 	 	 	 <= GEEF96
 	 	 	when 1010000100=> 
 	 	 	 	 <= GFG0CG
 	 	 	when 1010000101=> 
 	 	 	 	 <= GBC231
 	 	 	when 1010000110=> 
 	 	 	 	 <= G89D00
 	 	 	when 1010000111=> 
 	 	 	 	 <= GCCG4F
 	 	 	when 1010001000=> 
 	 	 	 	 <= GFF5B7
 	 	 	when 1010001001=> 
 	 	 	 	 <= GBC12F
 	 	 	when 1010001010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010001011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010001100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010001101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010001110=> 
 	 	 	 	 <= GDE178
 	 	 	when 1010001111=> 
 	 	 	 	 <= GBC230
 	 	 	when 1010010000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010010001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010010010=> 
 	 	 	 	 <= GCC83G
 	 	 	when 1010010011=> 
 	 	 	 	 <= GEEB8E
 	 	 	when 1010010100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010010101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010010110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010010111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010011000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010011001=> 
 	 	 	 	 <= G89D00
 	 	 	when 1010011010=> 
 	 	 	 	 <= GEEF97
 	 	 	when 1010011011=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1010011100=> 
 	 	 	 	 <= G9B412
 	 	 	when 1010011101=> 
 	 	 	 	 <= G9B311
 	 	 	when 1010011110=> 
 	 	 	 	 <= GFGFGE
 	 	 	when 1010100001=> 
 	 	 	 	 <= GFG5F5
 	 	 	when 1010100010=> 
 	 	 	 	 <= G99E01
 	 	 	when 1010100011=> 
 	 	 	 	 <= GBC73D
 	 	 	when 1010100100=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1010100101=> 
 	 	 	 	 <= GFFGCE
 	 	 	when 1010100110=> 
 	 	 	 	 <= GEF19E
 	 	 	when 1010100111=> 
 	 	 	 	 <= GDE47F
 	 	 	when 1010101000=> 
 	 	 	 	 <= G9B009
 	 	 	when 1010101001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010101010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010101011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010101100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010101101=> 
 	 	 	 	 <= G99D00
 	 	 	when 1010101110=> 
 	 	 	 	 <= GFF4B4
 	 	 	when 1010101111=> 
 	 	 	 	 <= G9B007
 	 	 	when 1010110000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010110001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010110010=> 
 	 	 	 	 <= G99D00
 	 	 	when 1010110011=> 
 	 	 	 	 <= GDE077
 	 	 	when 1010110100=> 
 	 	 	 	 <= GCD257
 	 	 	when 1010110101=> 
 	 	 	 	 <= G99D00
 	 	 	when 1010110110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010110111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010111000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1010111001=> 
 	 	 	 	 <= GBC334
 	 	 	when 1010111010=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1010111011=> 
 	 	 	 	 <= GEE683
 	 	 	when 1010111100=> 
 	 	 	 	 <= G99D00
 	 	 	when 1010111101=> 
 	 	 	 	 <= GCD870
 	 	 	when 1010111110=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1011000010=> 
 	 	 	 	 <= GCCF58
 	 	 	when 1011000011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011000100=> 
 	 	 	 	 <= GEEG99
 	 	 	when 1011000101=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1011000110=> 
 	 	 	 	 <= GEF19E
 	 	 	when 1011000111=> 
 	 	 	 	 <= G99D00
 	 	 	when 1011001000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011001001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011001010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011001011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011001100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011001101=> 
 	 	 	 	 <= G99G06
 	 	 	when 1011001110=> 
 	 	 	 	 <= GFF4B5
 	 	 	when 1011001111=> 
 	 	 	 	 <= G99D00
 	 	 	when 1011010000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011010001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011010010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011010011=> 
 	 	 	 	 <= G99G06
 	 	 	when 1011010100=> 
 	 	 	 	 <= GFF3B3
 	 	 	when 1011010101=> 
 	 	 	 	 <= GBBD24
 	 	 	when 1011010110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011010111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011011000=> 
 	 	 	 	 <= G9B009
 	 	 	when 1011011001=> 
 	 	 	 	 <= GFF7BC
 	 	 	when 1011011010=> 
 	 	 	 	 <= GFFGCF
 	 	 	when 1011011011=> 
 	 	 	 	 <= G9B81C
 	 	 	when 1011011100=> 
 	 	 	 	 <= G99F03
 	 	 	when 1011011101=> 
 	 	 	 	 <= GFG4F4
 	 	 	when 1011100010=> 
 	 	 	 	 <= GFG4F2
 	 	 	when 1011100011=> 
 	 	 	 	 <= G99G06
 	 	 	when 1011100100=> 
 	 	 	 	 <= G9B91D
 	 	 	when 1011100101=> 
 	 	 	 	 <= GFFFCC
 	 	 	when 1011100110=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1011100111=> 
 	 	 	 	 <= G9BC21
 	 	 	when 1011101000=> 
 	 	 	 	 <= G99D00
 	 	 	when 1011101001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011101010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011101011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011101100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011101101=> 
 	 	 	 	 <= GBC12G
 	 	 	when 1011101110=> 
 	 	 	 	 <= GDE27B
 	 	 	when 1011101111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011110000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011110001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011110010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011110011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011110100=> 
 	 	 	 	 <= GBBC21
 	 	 	when 1011110101=> 
 	 	 	 	 <= GFF4B5
 	 	 	when 1011110110=> 
 	 	 	 	 <= G9B007
 	 	 	when 1011110111=> 
 	 	 	 	 <= G99F03
 	 	 	when 1011111000=> 
 	 	 	 	 <= GEEB8F
 	 	 	when 1011111001=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1011111010=> 
 	 	 	 	 <= GCD45C
 	 	 	when 1011111011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1011111100=> 
 	 	 	 	 <= GCD973
 	 	 	when 1011111101=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1100000011=> 
 	 	 	 	 <= GDE594
 	 	 	when 1100000100=> 
 	 	 	 	 <= G89D00
 	 	 	when 1100000101=> 
 	 	 	 	 <= GCC73F
 	 	 	when 1100000110=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1100000111=> 
 	 	 	 	 <= GFFCC3
 	 	 	when 1100001000=> 
 	 	 	 	 <= GBBE26
 	 	 	when 1100001001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100001010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100001011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100001100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100001101=> 
 	 	 	 	 <= GCD45C
 	 	 	when 1100001110=> 
 	 	 	 	 <= GCCG4F
 	 	 	when 1100001111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100010000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100010001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100010010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100010011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100010100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100010101=> 
 	 	 	 	 <= GCD153
 	 	 	when 1100010110=> 
 	 	 	 	 <= GEF19F
 	 	 	when 1100010111=> 
 	 	 	 	 <= GEF2B0
 	 	 	when 1100011000=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1100011001=> 
 	 	 	 	 <= GEE582
 	 	 	when 1100011010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100011011=> 
 	 	 	 	 <= G9BB23
 	 	 	when 1100011100=> 
 	 	 	 	 <= GFGDG7
 	 	 	when 1100100011=> 
 	 	 	 	 <= GGGFGF
 	 	 	when 1100100100=> 
 	 	 	 	 <= GCD05C
 	 	 	when 1100100101=> 
 	 	 	 	 <= G99D00
 	 	 	when 1100100110=> 
 	 	 	 	 <= GCCC46
 	 	 	when 1100100111=> 
 	 	 	 	 <= GFG0CG
 	 	 	when 1100101000=> 
 	 	 	 	 <= GFFGCE
 	 	 	when 1100101001=> 
 	 	 	 	 <= GCD55D
 	 	 	when 1100101010=> 
 	 	 	 	 <= G99F03
 	 	 	when 1100101011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100101100=> 
 	 	 	 	 <= G99D00
 	 	 	when 1100101101=> 
 	 	 	 	 <= GEE787
 	 	 	when 1100101110=> 
 	 	 	 	 <= GBBC22
 	 	 	when 1100101111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100110000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100110001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100110010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100110011=> 
 	 	 	 	 <= G99E00
 	 	 	when 1100110100=> 
 	 	 	 	 <= G99D00
 	 	 	when 1100110101=> 
 	 	 	 	 <= GCCG50
 	 	 	when 1100110110=> 
 	 	 	 	 <= GGG0D1
 	 	 	when 1100110111=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 1100111000=> 
 	 	 	 	 <= GEE582
 	 	 	when 1100111001=> 
 	 	 	 	 <= G99F02
 	 	 	when 1100111010=> 
 	 	 	 	 <= G9B10D
 	 	 	when 1100111011=> 
 	 	 	 	 <= GFG0E9
 	 	 	when 1101000100=> 
 	 	 	 	 <= GFGEGC
 	 	 	when 1101000101=> 
 	 	 	 	 <= GBCC4F
 	 	 	when 1101000110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1101000111=> 
 	 	 	 	 <= GBC02D
 	 	 	when 1101001000=> 
 	 	 	 	 <= GFF8BE
 	 	 	when 1101001001=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1101001010=> 
 	 	 	 	 <= GFF9BG
 	 	 	when 1101001011=> 
 	 	 	 	 <= GCD55D
 	 	 	when 1101001100=> 
 	 	 	 	 <= GBC230
 	 	 	when 1101001101=> 
 	 	 	 	 <= GFFDC6
 	 	 	when 1101001110=> 
 	 	 	 	 <= G9B719
 	 	 	when 1101001111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1101010000=> 
 	 	 	 	 <= G99E00
 	 	 	when 1101010001=> 
 	 	 	 	 <= G99E00
 	 	 	when 1101010010=> 
 	 	 	 	 <= G9B008
 	 	 	when 1101010011=> 
 	 	 	 	 <= GCC942
 	 	 	when 1101010100=> 
 	 	 	 	 <= GEEE95
 	 	 	when 1101010101=> 
 	 	 	 	 <= GFG0D1
 	 	 	when 1101010110=> 
 	 	 	 	 <= GFFGCF
 	 	 	when 1101010111=> 
 	 	 	 	 <= GCD45C
 	 	 	when 1101011000=> 
 	 	 	 	 <= G89E00
 	 	 	when 1101011001=> 
 	 	 	 	 <= G9B10D
 	 	 	when 1101011010=> 
 	 	 	 	 <= GEFCDC
 	 	 	when 1101100101=> 
 	 	 	 	 <= GFGFGE
 	 	 	when 1101100110=> 
 	 	 	 	 <= GCD871
 	 	 	when 1101100111=> 
 	 	 	 	 <= G99D00
 	 	 	when 1101101000=> 
 	 	 	 	 <= G99G06
 	 	 	when 1101101001=> 
 	 	 	 	 <= GDD762
 	 	 	when 1101101010=> 
 	 	 	 	 <= GFFDC7
 	 	 	when 1101101011=> 
 	 	 	 	 <= GFG1D1
 	 	 	when 1101101100=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1101101101=> 
 	 	 	 	 <= GGG1D1
 	 	 	when 1101101110=> 
 	 	 	 	 <= GFFFCC
 	 	 	when 1101101111=> 
 	 	 	 	 <= GEEF96
 	 	 	when 1101110000=> 
 	 	 	 	 <= GEEF96
 	 	 	when 1101110001=> 
 	 	 	 	 <= GFF6B7
 	 	 	when 1101110010=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1101110011=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1101110100=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1101110101=> 
 	 	 	 	 <= GEE785
 	 	 	when 1101110110=> 
 	 	 	 	 <= G9B91D
 	 	 	when 1101110111=> 
 	 	 	 	 <= G99D00
 	 	 	when 1101111000=> 
 	 	 	 	 <= G9BB24
 	 	 	when 1101111001=> 
 	 	 	 	 <= GFG0EB
 	 	 	when 1110000110=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1110000111=> 
 	 	 	 	 <= GEF5CC
 	 	 	when 1110001000=> 
 	 	 	 	 <= G9B920
 	 	 	when 1110001001=> 
 	 	 	 	 <= G99D00
 	 	 	when 1110001010=> 
 	 	 	 	 <= G99G05
 	 	 	when 1110001011=> 
 	 	 	 	 <= GCC942
 	 	 	when 1110001100=> 
 	 	 	 	 <= GDE37D
 	 	 	when 1110001101=> 
 	 	 	 	 <= GFF5B6
 	 	 	when 1110001110=> 
 	 	 	 	 <= GFFGCF
 	 	 	when 1110001111=> 
 	 	 	 	 <= GGG0D1
 	 	 	when 1110010000=> 
 	 	 	 	 <= GFG0D0
 	 	 	when 1110010001=> 
 	 	 	 	 <= GFFBC1
 	 	 	when 1110010010=> 
 	 	 	 	 <= GEEB8E
 	 	 	when 1110010011=> 
 	 	 	 	 <= GCD358
 	 	 	when 1110010100=> 
 	 	 	 	 <= G9B614
 	 	 	when 1110010101=> 
 	 	 	 	 <= G99E00
 	 	 	when 1110010110=> 
 	 	 	 	 <= G99F02
 	 	 	when 1110010111=> 
 	 	 	 	 <= GCD770
 	 	 	when 1110011000=> 
 	 	 	 	 <= GFGCG7
 	 	 	when 1110101000=> 
 	 	 	 	 <= GFGEGD
 	 	 	when 1110101001=> 
 	 	 	 	 <= GDEBB0
 	 	 	when 1110101010=> 
 	 	 	 	 <= GBBG30
 	 	 	when 1110101011=> 
 	 	 	 	 <= G99D00
 	 	 	when 1110101100=> 
 	 	 	 	 <= G99E00
 	 	 	when 1110101101=> 
 	 	 	 	 <= G89D00
 	 	 	when 1110101110=> 
 	 	 	 	 <= G99E00
 	 	 	when 1110101111=> 
 	 	 	 	 <= G99E00
 	 	 	when 1110110000=> 
 	 	 	 	 <= G99D00
 	 	 	when 1110110001=> 
 	 	 	 	 <= G89D00
 	 	 	when 1110110010=> 
 	 	 	 	 <= G99E00
 	 	 	when 1110110011=> 
 	 	 	 	 <= G89D00
 	 	 	when 1110110100=> 
 	 	 	 	 <= G9B10D
 	 	 	when 1110110101=> 
 	 	 	 	 <= GCD56B
 	 	 	when 1110110110=> 
 	 	 	 	 <= GFG3F0
 	 	 	when 1110110111=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1111001010=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1111001011=> 
 	 	 	 	 <= GFG4F4
 	 	 	when 1111001100=> 
 	 	 	 	 <= GDEB9G
 	 	 	when 1111001101=> 
 	 	 	 	 <= GCD76E
 	 	 	when 1111001110=> 
 	 	 	 	 <= GBCB4F
 	 	 	when 1111001111=> 
 	 	 	 	 <= GBC540
 	 	 	when 1111010000=> 
 	 	 	 	 <= GBC847
 	 	 	when 1111010001=> 
 	 	 	 	 <= GCD05D
 	 	 	when 1111010010=> 
 	 	 	 	 <= GDE085
 	 	 	when 1111010011=> 
 	 	 	 	 <= GEF7D2
 	 	 	when 1111010100=> 
 	 	 	 	 <= GFGEGD
 	 	 	when 1111010101=> 
 	 	 	 	 <= GFGFGF 
 	 	 end case; 
     	 end if;  
     end process; 
 address <= row & col; 
 end;