library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity CHERRYROM is
  port(
	  row : in std_logic_vector(4 downto 0);
	  col : in std_logic_vector(4 downto 0);
	  fruit_color : in std_logic_vector(5 downto 0);
	  clk : in std_logic;
	  color : out std_logic_vector(5 downto 0)
  );
end CHERRYROM;

architecture synth of CHERRYROM is 
signal address : std_logic_vector(9 downto 0);
begin
	process(clk) is
	begin
		if rising_edge(clk) then
			case address is 

 	 	 	when 0000001110=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000001111=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000010000=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0000101010=> 
 	 	 	 	 <= G9FGFG
 	 	 	when 0000101011=> 
 	 	 	 	 <= F3B9B9
 	 	 	when 0000101100=> 
 	 	 	 	 <= E16G6G
 	 	 	when 0000101101=> 
 	 	 	 	 <= D44444
 	 	 	when 0000101110=> 
 	 	 	 	 <= CC2929
 	 	 	when 0000101111=> 
 	 	 	 	 <= C81G20
 	 	 	when 0000110000=> 
 	 	 	 	 <= C92121
 	 	 	when 0000110001=> 
 	 	 	 	 <= CF3434
 	 	 	when 0000110010=> 
 	 	 	 	 <= D95454
 	 	 	when 0000110011=> 
 	 	 	 	 <= E88686
 	 	 	when 0000110100=> 
 	 	 	 	 <= FED8D8
 	 	 	when 0000110101=> 
 	 	 	 	 <= GFGEGE
 	 	 	when 0001001000=> 
 	 	 	 	 <= FFD9D9
 	 	 	when 0001001001=> 
 	 	 	 	 <= DB5959
 	 	 	when 0001001010=> 
 	 	 	 	 <= C51616
 	 	 	when 0001001011=> 
 	 	 	 	 <= C51515
 	 	 	when 0001001100=> 
 	 	 	 	 <= C51515
 	 	 	when 0001001101=> 
 	 	 	 	 <= C51515
 	 	 	when 0001001110=> 
 	 	 	 	 <= C51515
 	 	 	when 0001001111=> 
 	 	 	 	 <= C51515
 	 	 	when 0001010000=> 
 	 	 	 	 <= C51515
 	 	 	when 0001010001=> 
 	 	 	 	 <= C51515
 	 	 	when 0001010010=> 
 	 	 	 	 <= C51515
 	 	 	when 0001010011=> 
 	 	 	 	 <= C51515
 	 	 	when 0001010100=> 
 	 	 	 	 <= C51515
 	 	 	when 0001010101=> 
 	 	 	 	 <= CC2828
 	 	 	when 0001010110=> 
 	 	 	 	 <= E98989
 	 	 	when 0001010111=> 
 	 	 	 	 <= GBG1G1
 	 	 	when 0001100110=> 
 	 	 	 	 <= G7F6F6
 	 	 	when 0001100111=> 
 	 	 	 	 <= DB5757
 	 	 	when 0001101000=> 
 	 	 	 	 <= C51415
 	 	 	when 0001101001=> 
 	 	 	 	 <= C51515
 	 	 	when 0001101010=> 
 	 	 	 	 <= C51515
 	 	 	when 0001101011=> 
 	 	 	 	 <= C51515
 	 	 	when 0001101100=> 
 	 	 	 	 <= C51515
 	 	 	when 0001101101=> 
 	 	 	 	 <= C51515
 	 	 	when 0001101110=> 
 	 	 	 	 <= C51515
 	 	 	when 0001101111=> 
 	 	 	 	 <= C51515
 	 	 	when 0001110000=> 
 	 	 	 	 <= C51515
 	 	 	when 0001110001=> 
 	 	 	 	 <= C51515
 	 	 	when 0001110010=> 
 	 	 	 	 <= C51515
 	 	 	when 0001110011=> 
 	 	 	 	 <= C51515
 	 	 	when 0001110100=> 
 	 	 	 	 <= C51515
 	 	 	when 0001110101=> 
 	 	 	 	 <= C51515
 	 	 	when 0001110110=> 
 	 	 	 	 <= C51515
 	 	 	when 0001110111=> 
 	 	 	 	 <= C82020
 	 	 	when 0001111000=> 
 	 	 	 	 <= EG9C9C
 	 	 	when 0001111001=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0010000100=> 
 	 	 	 	 <= GFGFGG
 	 	 	when 0010000101=> 
 	 	 	 	 <= F8C7C7
 	 	 	when 0010000110=> 
 	 	 	 	 <= C81G1G
 	 	 	when 0010000111=> 
 	 	 	 	 <= C51515
 	 	 	when 0010001000=> 
 	 	 	 	 <= C51515
 	 	 	when 0010001001=> 
 	 	 	 	 <= C51415
 	 	 	when 0010001010=> 
 	 	 	 	 <= C41414
 	 	 	when 0010001011=> 
 	 	 	 	 <= C51515
 	 	 	when 0010001100=> 
 	 	 	 	 <= C51515
 	 	 	when 0010001101=> 
 	 	 	 	 <= C51515
 	 	 	when 0010001110=> 
 	 	 	 	 <= C51515
 	 	 	when 0010001111=> 
 	 	 	 	 <= C51515
 	 	 	when 0010010000=> 
 	 	 	 	 <= C51515
 	 	 	when 0010010001=> 
 	 	 	 	 <= C51515
 	 	 	when 0010010010=> 
 	 	 	 	 <= C51515
 	 	 	when 0010010011=> 
 	 	 	 	 <= C51515
 	 	 	when 0010010100=> 
 	 	 	 	 <= C51515
 	 	 	when 0010010101=> 
 	 	 	 	 <= C51515
 	 	 	when 0010010110=> 
 	 	 	 	 <= C51515
 	 	 	when 0010010111=> 
 	 	 	 	 <= C51515
 	 	 	when 0010011000=> 
 	 	 	 	 <= C51515
 	 	 	when 0010011001=> 
 	 	 	 	 <= D74G50
 	 	 	when 0010011010=> 
 	 	 	 	 <= GBG0G0
 	 	 	when 0010100011=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0010100100=> 
 	 	 	 	 <= F09G9G
 	 	 	when 0010100101=> 
 	 	 	 	 <= C51515
 	 	 	when 0010100110=> 
 	 	 	 	 <= C51515
 	 	 	when 0010100111=> 
 	 	 	 	 <= C51515
 	 	 	when 0010101000=> 
 	 	 	 	 <= BG1414
 	 	 	when 0010101001=> 
 	 	 	 	 <= 790D0D
 	 	 	when 0010101010=> 
 	 	 	 	 <= 850F0F
 	 	 	when 0010101011=> 
 	 	 	 	 <= C51515
 	 	 	when 0010101100=> 
 	 	 	 	 <= C51515
 	 	 	when 0010101101=> 
 	 	 	 	 <= C51515
 	 	 	when 0010101110=> 
 	 	 	 	 <= C51515
 	 	 	when 0010101111=> 
 	 	 	 	 <= C51515
 	 	 	when 0010110000=> 
 	 	 	 	 <= C51515
 	 	 	when 0010110001=> 
 	 	 	 	 <= C51515
 	 	 	when 0010110010=> 
 	 	 	 	 <= C51515
 	 	 	when 0010110011=> 
 	 	 	 	 <= C51515
 	 	 	when 0010110100=> 
 	 	 	 	 <= C51515
 	 	 	when 0010110101=> 
 	 	 	 	 <= C51515
 	 	 	when 0010110110=> 
 	 	 	 	 <= C51515
 	 	 	when 0010110111=> 
 	 	 	 	 <= C51515
 	 	 	when 0010111000=> 
 	 	 	 	 <= C51515
 	 	 	when 0010111001=> 
 	 	 	 	 <= C51515
 	 	 	when 0010111010=> 
 	 	 	 	 <= CF3434
 	 	 	when 0010111011=> 
 	 	 	 	 <= G7F8F8
 	 	 	when 0011000011=> 
 	 	 	 	 <= F5BEBE
 	 	 	when 0011000100=> 
 	 	 	 	 <= C51515
 	 	 	when 0011000101=> 
 	 	 	 	 <= C51515
 	 	 	when 0011000110=> 
 	 	 	 	 <= C51515
 	 	 	when 0011000111=> 
 	 	 	 	 <= C21414
 	 	 	when 0011001000=> 
 	 	 	 	 <= 790D0D
 	 	 	when 0011001001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0011001010=> 
 	 	 	 	 <= 770D0D
 	 	 	when 0011001011=> 
 	 	 	 	 <= C51515
 	 	 	when 0011001100=> 
 	 	 	 	 <= C51515
 	 	 	when 0011001101=> 
 	 	 	 	 <= C51515
 	 	 	when 0011001110=> 
 	 	 	 	 <= C51515
 	 	 	when 0011001111=> 
 	 	 	 	 <= C51515
 	 	 	when 0011010000=> 
 	 	 	 	 <= C51515
 	 	 	when 0011010001=> 
 	 	 	 	 <= C51515
 	 	 	when 0011010010=> 
 	 	 	 	 <= C51515
 	 	 	when 0011010011=> 
 	 	 	 	 <= C51515
 	 	 	when 0011010100=> 
 	 	 	 	 <= C51515
 	 	 	when 0011010101=> 
 	 	 	 	 <= C51515
 	 	 	when 0011010110=> 
 	 	 	 	 <= C51515
 	 	 	when 0011010111=> 
 	 	 	 	 <= C51515
 	 	 	when 0011011000=> 
 	 	 	 	 <= C51515
 	 	 	when 0011011001=> 
 	 	 	 	 <= C51515
 	 	 	when 0011011010=> 
 	 	 	 	 <= C51515
 	 	 	when 0011011011=> 
 	 	 	 	 <= CG3636
 	 	 	when 0011011100=> 
 	 	 	 	 <= GCG3G3
 	 	 	when 0011100010=> 
 	 	 	 	 <= G2EBEB
 	 	 	when 0011100011=> 
 	 	 	 	 <= 8G1414
 	 	 	when 0011100100=> 
 	 	 	 	 <= 790D0D
 	 	 	when 0011100101=> 
 	 	 	 	 <= 860F0F
 	 	 	when 0011100110=> 
 	 	 	 	 <= 921010
 	 	 	when 0011100111=> 
 	 	 	 	 <= 710C0C
 	 	 	when 0011101000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0011101001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0011101010=> 
 	 	 	 	 <= 991111
 	 	 	when 0011101011=> 
 	 	 	 	 <= C51515
 	 	 	when 0011101100=> 
 	 	 	 	 <= C51515
 	 	 	when 0011101101=> 
 	 	 	 	 <= C51515
 	 	 	when 0011101110=> 
 	 	 	 	 <= C51515
 	 	 	when 0011101111=> 
 	 	 	 	 <= C51515
 	 	 	when 0011110000=> 
 	 	 	 	 <= C51515
 	 	 	when 0011110001=> 
 	 	 	 	 <= C51515
 	 	 	when 0011110010=> 
 	 	 	 	 <= C51515
 	 	 	when 0011110011=> 
 	 	 	 	 <= C51515
 	 	 	when 0011110100=> 
 	 	 	 	 <= C51515
 	 	 	when 0011110101=> 
 	 	 	 	 <= C51515
 	 	 	when 0011110110=> 
 	 	 	 	 <= C51515
 	 	 	when 0011110111=> 
 	 	 	 	 <= C51515
 	 	 	when 0011111000=> 
 	 	 	 	 <= C51515
 	 	 	when 0011111001=> 
 	 	 	 	 <= C51515
 	 	 	when 0011111010=> 
 	 	 	 	 <= C51515
 	 	 	when 0011111011=> 
 	 	 	 	 <= C51515
 	 	 	when 0011111100=> 
 	 	 	 	 <= DB5959
 	 	 	when 0011111101=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0100000001=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 0100000010=> 
 	 	 	 	 <= 8G3C3C
 	 	 	when 0100000011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0100000100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0100000101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0100000110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0100000111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0100001000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0100001001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0100001010=> 
 	 	 	 	 <= B61212
 	 	 	when 0100001011=> 
 	 	 	 	 <= C51515
 	 	 	when 0100001100=> 
 	 	 	 	 <= C51515
 	 	 	when 0100001101=> 
 	 	 	 	 <= C51515
 	 	 	when 0100001110=> 
 	 	 	 	 <= C51515
 	 	 	when 0100001111=> 
 	 	 	 	 <= C51515
 	 	 	when 0100010000=> 
 	 	 	 	 <= C51515
 	 	 	when 0100010001=> 
 	 	 	 	 <= C51515
 	 	 	when 0100010010=> 
 	 	 	 	 <= C51515
 	 	 	when 0100010011=> 
 	 	 	 	 <= C51515
 	 	 	when 0100010100=> 
 	 	 	 	 <= C51515
 	 	 	when 0100010101=> 
 	 	 	 	 <= C51515
 	 	 	when 0100010110=> 
 	 	 	 	 <= C51515
 	 	 	when 0100010111=> 
 	 	 	 	 <= C51515
 	 	 	when 0100011000=> 
 	 	 	 	 <= C51515
 	 	 	when 0100011001=> 
 	 	 	 	 <= C51515
 	 	 	when 0100011010=> 
 	 	 	 	 <= C51515
 	 	 	when 0100011011=> 
 	 	 	 	 <= C51515
 	 	 	when 0100011100=> 
 	 	 	 	 <= C41414
 	 	 	when 0100011101=> 
 	 	 	 	 <= F5BEBE
 	 	 	when 0100100001=> 
 	 	 	 	 <= D29E9E
 	 	 	when 0100100010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0100100011=> 
 	 	 	 	 <= 6D0B0B
 	 	 	when 0100100100=> 
 	 	 	 	 <= B31212
 	 	 	when 0100100101=> 
 	 	 	 	 <= 750C0C
 	 	 	when 0100100110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0100100111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0100101000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0100101001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0100101010=> 
 	 	 	 	 <= BB1313
 	 	 	when 0100101011=> 
 	 	 	 	 <= C51515
 	 	 	when 0100101100=> 
 	 	 	 	 <= C51515
 	 	 	when 0100101101=> 
 	 	 	 	 <= C51515
 	 	 	when 0100101110=> 
 	 	 	 	 <= C51515
 	 	 	when 0100101111=> 
 	 	 	 	 <= C51515
 	 	 	when 0100110000=> 
 	 	 	 	 <= C51515
 	 	 	when 0100110001=> 
 	 	 	 	 <= C51515
 	 	 	when 0100110010=> 
 	 	 	 	 <= C51515
 	 	 	when 0100110011=> 
 	 	 	 	 <= C51515
 	 	 	when 0100110100=> 
 	 	 	 	 <= C51515
 	 	 	when 0100110101=> 
 	 	 	 	 <= C51515
 	 	 	when 0100110110=> 
 	 	 	 	 <= C51515
 	 	 	when 0100110111=> 
 	 	 	 	 <= C51515
 	 	 	when 0100111000=> 
 	 	 	 	 <= C51515
 	 	 	when 0100111001=> 
 	 	 	 	 <= C51515
 	 	 	when 0100111010=> 
 	 	 	 	 <= C51515
 	 	 	when 0100111011=> 
 	 	 	 	 <= C51515
 	 	 	when 0100111100=> 
 	 	 	 	 <= C51515
 	 	 	when 0100111101=> 
 	 	 	 	 <= CD2D2D
 	 	 	when 0100111110=> 
 	 	 	 	 <= GEGCGC
 	 	 	when 0101000000=> 
 	 	 	 	 <= GFGEGE
 	 	 	when 0101000001=> 
 	 	 	 	 <= 782424
 	 	 	when 0101000010=> 
 	 	 	 	 <= 690B0B
 	 	 	when 0101000011=> 
 	 	 	 	 <= B51212
 	 	 	when 0101000100=> 
 	 	 	 	 <= C51515
 	 	 	when 0101000101=> 
 	 	 	 	 <= BD1313
 	 	 	when 0101000110=> 
 	 	 	 	 <= 6D0B0B
 	 	 	when 0101000111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0101001000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0101001001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0101001010=> 
 	 	 	 	 <= B81313
 	 	 	when 0101001011=> 
 	 	 	 	 <= C51515
 	 	 	when 0101001100=> 
 	 	 	 	 <= C51515
 	 	 	when 0101001101=> 
 	 	 	 	 <= C51515
 	 	 	when 0101001110=> 
 	 	 	 	 <= C51515
 	 	 	when 0101001111=> 
 	 	 	 	 <= C51515
 	 	 	when 0101010000=> 
 	 	 	 	 <= C51515
 	 	 	when 0101010001=> 
 	 	 	 	 <= C51515
 	 	 	when 0101010010=> 
 	 	 	 	 <= C51515
 	 	 	when 0101010011=> 
 	 	 	 	 <= C51515
 	 	 	when 0101010100=> 
 	 	 	 	 <= C51515
 	 	 	when 0101010101=> 
 	 	 	 	 <= C51515
 	 	 	when 0101010110=> 
 	 	 	 	 <= C51515
 	 	 	when 0101010111=> 
 	 	 	 	 <= C51515
 	 	 	when 0101011000=> 
 	 	 	 	 <= C51515
 	 	 	when 0101011001=> 
 	 	 	 	 <= C51515
 	 	 	when 0101011010=> 
 	 	 	 	 <= C51515
 	 	 	when 0101011011=> 
 	 	 	 	 <= C51515
 	 	 	when 0101011100=> 
 	 	 	 	 <= C51515
 	 	 	when 0101011101=> 
 	 	 	 	 <= C51515
 	 	 	when 0101011110=> 
 	 	 	 	 <= F4BDBD
 	 	 	when 0101100000=> 
 	 	 	 	 <= FBE2E2
 	 	 	when 0101100001=> 
 	 	 	 	 <= 700C0C
 	 	 	when 0101100010=> 
 	 	 	 	 <= 910G0G
 	 	 	when 0101100011=> 
 	 	 	 	 <= C51415
 	 	 	when 0101100100=> 
 	 	 	 	 <= C41414
 	 	 	when 0101100101=> 
 	 	 	 	 <= C51515
 	 	 	when 0101100110=> 
 	 	 	 	 <= 951010
 	 	 	when 0101100111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0101101000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0101101001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0101101010=> 
 	 	 	 	 <= 9F1111
 	 	 	when 0101101011=> 
 	 	 	 	 <= C51515
 	 	 	when 0101101100=> 
 	 	 	 	 <= C51515
 	 	 	when 0101101101=> 
 	 	 	 	 <= B61212
 	 	 	when 0101101110=> 
 	 	 	 	 <= 8F0G0G
 	 	 	when 0101101111=> 
 	 	 	 	 <= 92100G
 	 	 	when 0101110000=> 
 	 	 	 	 <= C41414
 	 	 	when 0101110001=> 
 	 	 	 	 <= C51515
 	 	 	when 0101110010=> 
 	 	 	 	 <= C51515
 	 	 	when 0101110011=> 
 	 	 	 	 <= C51515
 	 	 	when 0101110100=> 
 	 	 	 	 <= C51515
 	 	 	when 0101110101=> 
 	 	 	 	 <= C51515
 	 	 	when 0101110110=> 
 	 	 	 	 <= C51515
 	 	 	when 0101110111=> 
 	 	 	 	 <= C51515
 	 	 	when 0101111000=> 
 	 	 	 	 <= C51515
 	 	 	when 0101111001=> 
 	 	 	 	 <= C51515
 	 	 	when 0101111010=> 
 	 	 	 	 <= C51515
 	 	 	when 0101111011=> 
 	 	 	 	 <= C51515
 	 	 	when 0101111100=> 
 	 	 	 	 <= C51515
 	 	 	when 0101111101=> 
 	 	 	 	 <= C51515
 	 	 	when 0101111110=> 
 	 	 	 	 <= D85151
 	 	 	when 0110000000=> 
 	 	 	 	 <= EE9595
 	 	 	when 0110000001=> 
 	 	 	 	 <= C51414
 	 	 	when 0110000010=> 
 	 	 	 	 <= C41414
 	 	 	when 0110000011=> 
 	 	 	 	 <= 8B0F0F
 	 	 	when 0110000100=> 
 	 	 	 	 <= 880F0F
 	 	 	when 0110000101=> 
 	 	 	 	 <= C41414
 	 	 	when 0110000110=> 
 	 	 	 	 <= C41414
 	 	 	when 0110000111=> 
 	 	 	 	 <= 6E0B0B
 	 	 	when 0110001000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0110001001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0110001010=> 
 	 	 	 	 <= 9B1111
 	 	 	when 0110001011=> 
 	 	 	 	 <= C51515
 	 	 	when 0110001100=> 
 	 	 	 	 <= C51515
 	 	 	when 0110001101=> 
 	 	 	 	 <= 7B0D0D
 	 	 	when 0110001110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0110001111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0110010000=> 
 	 	 	 	 <= 9D1111
 	 	 	when 0110010001=> 
 	 	 	 	 <= C51515
 	 	 	when 0110010010=> 
 	 	 	 	 <= C51515
 	 	 	when 0110010011=> 
 	 	 	 	 <= C51515
 	 	 	when 0110010100=> 
 	 	 	 	 <= C51515
 	 	 	when 0110010101=> 
 	 	 	 	 <= C51515
 	 	 	when 0110010110=> 
 	 	 	 	 <= C51515
 	 	 	when 0110010111=> 
 	 	 	 	 <= C51515
 	 	 	when 0110011000=> 
 	 	 	 	 <= C51515
 	 	 	when 0110011001=> 
 	 	 	 	 <= C51515
 	 	 	when 0110011010=> 
 	 	 	 	 <= C51515
 	 	 	when 0110011011=> 
 	 	 	 	 <= C51515
 	 	 	when 0110011100=> 
 	 	 	 	 <= C41414
 	 	 	when 0110011101=> 
 	 	 	 	 <= C51414
 	 	 	when 0110011110=> 
 	 	 	 	 <= C61818
 	 	 	when 0110100000=> 
 	 	 	 	 <= DE6363
 	 	 	when 0110100001=> 
 	 	 	 	 <= C51515
 	 	 	when 0110100010=> 
 	 	 	 	 <= 9D1111
 	 	 	when 0110100011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0110100100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0110100101=> 
 	 	 	 	 <= B21212
 	 	 	when 0110100110=> 
 	 	 	 	 <= C51515
 	 	 	when 0110100111=> 
 	 	 	 	 <= 7G0E0E
 	 	 	when 0110101000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0110101001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0110101010=> 
 	 	 	 	 <= 981010
 	 	 	when 0110101011=> 
 	 	 	 	 <= C51515
 	 	 	when 0110101100=> 
 	 	 	 	 <= C51515
 	 	 	when 0110101101=> 
 	 	 	 	 <= 900G0G
 	 	 	when 0110101110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0110101111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0110110000=> 
 	 	 	 	 <= 971010
 	 	 	when 0110110001=> 
 	 	 	 	 <= C51515
 	 	 	when 0110110010=> 
 	 	 	 	 <= C51515
 	 	 	when 0110110011=> 
 	 	 	 	 <= C51515
 	 	 	when 0110110100=> 
 	 	 	 	 <= C51515
 	 	 	when 0110110101=> 
 	 	 	 	 <= C51515
 	 	 	when 0110110110=> 
 	 	 	 	 <= C51515
 	 	 	when 0110110111=> 
 	 	 	 	 <= C51515
 	 	 	when 0110111000=> 
 	 	 	 	 <= C51515
 	 	 	when 0110111001=> 
 	 	 	 	 <= C51515
 	 	 	when 0110111010=> 
 	 	 	 	 <= C51515
 	 	 	when 0110111011=> 
 	 	 	 	 <= C51515
 	 	 	when 0110111100=> 
 	 	 	 	 <= B11212
 	 	 	when 0110111101=> 
 	 	 	 	 <= 770D0D
 	 	 	when 0110111110=> 
 	 	 	 	 <= B51212
 	 	 	when 0111000000=> 
 	 	 	 	 <= D34444
 	 	 	when 0111000001=> 
 	 	 	 	 <= C51515
 	 	 	when 0111000010=> 
 	 	 	 	 <= 8C0G0G
 	 	 	when 0111000011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0111000100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0111000101=> 
 	 	 	 	 <= 8C0G0G
 	 	 	when 0111000110=> 
 	 	 	 	 <= C51515
 	 	 	when 0111000111=> 
 	 	 	 	 <= 8E0G0G
 	 	 	when 0111001000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0111001001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0111001010=> 
 	 	 	 	 <= 971110
 	 	 	when 0111001011=> 
 	 	 	 	 <= C51515
 	 	 	when 0111001100=> 
 	 	 	 	 <= C51515
 	 	 	when 0111001101=> 
 	 	 	 	 <= BB1313
 	 	 	when 0111001110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0111001111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0111010000=> 
 	 	 	 	 <= 910G0G
 	 	 	when 0111010001=> 
 	 	 	 	 <= C51515
 	 	 	when 0111010010=> 
 	 	 	 	 <= C51515
 	 	 	when 0111010011=> 
 	 	 	 	 <= C51515
 	 	 	when 0111010100=> 
 	 	 	 	 <= C51515
 	 	 	when 0111010101=> 
 	 	 	 	 <= C51515
 	 	 	when 0111010110=> 
 	 	 	 	 <= C51515
 	 	 	when 0111010111=> 
 	 	 	 	 <= C51515
 	 	 	when 0111011000=> 
 	 	 	 	 <= C51515
 	 	 	when 0111011001=> 
 	 	 	 	 <= C51515
 	 	 	when 0111011010=> 
 	 	 	 	 <= C51515
 	 	 	when 0111011011=> 
 	 	 	 	 <= BG1414
 	 	 	when 0111011100=> 
 	 	 	 	 <= 6G0C0C
 	 	 	when 0111011101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0111011110=> 
 	 	 	 	 <= 8E0G0G
 	 	 	when 0111100000=> 
 	 	 	 	 <= CG3434
 	 	 	when 0111100001=> 
 	 	 	 	 <= C51515
 	 	 	when 0111100010=> 
 	 	 	 	 <= 820E0E
 	 	 	when 0111100011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0111100100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0111100101=> 
 	 	 	 	 <= 6B0B0B
 	 	 	when 0111100110=> 
 	 	 	 	 <= C21414
 	 	 	when 0111100111=> 
 	 	 	 	 <= 921010
 	 	 	when 0111101000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0111101001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0111101010=> 
 	 	 	 	 <= 971010
 	 	 	when 0111101011=> 
 	 	 	 	 <= C51515
 	 	 	when 0111101100=> 
 	 	 	 	 <= C51515
 	 	 	when 0111101101=> 
 	 	 	 	 <= C41414
 	 	 	when 0111101110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0111101111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0111110000=> 
 	 	 	 	 <= 880F0F
 	 	 	when 0111110001=> 
 	 	 	 	 <= C51515
 	 	 	when 0111110010=> 
 	 	 	 	 <= C51515
 	 	 	when 0111110011=> 
 	 	 	 	 <= C51515
 	 	 	when 0111110100=> 
 	 	 	 	 <= C51515
 	 	 	when 0111110101=> 
 	 	 	 	 <= C51515
 	 	 	when 0111110110=> 
 	 	 	 	 <= C51515
 	 	 	when 0111110111=> 
 	 	 	 	 <= C51515
 	 	 	when 0111111000=> 
 	 	 	 	 <= C51515
 	 	 	when 0111111001=> 
 	 	 	 	 <= C51515
 	 	 	when 0111111010=> 
 	 	 	 	 <= C41414
 	 	 	when 0111111011=> 
 	 	 	 	 <= 7B0D0D
 	 	 	when 0111111100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0111111101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 0111111110=> 
 	 	 	 	 <= 8E0G0G
 	 	 	when 1000000000=> 
 	 	 	 	 <= D03939
 	 	 	when 1000000001=> 
 	 	 	 	 <= C51515
 	 	 	when 1000000010=> 
 	 	 	 	 <= 840F0F
 	 	 	when 1000000011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1000000100=> 
 	 	 	 	 <= 690B0B
 	 	 	when 1000000101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1000000110=> 
 	 	 	 	 <= B41212
 	 	 	when 1000000111=> 
 	 	 	 	 <= 8B0F0F
 	 	 	when 1000001000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1000001001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1000001010=> 
 	 	 	 	 <= 951010
 	 	 	when 1000001011=> 
 	 	 	 	 <= C51515
 	 	 	when 1000001100=> 
 	 	 	 	 <= C51515
 	 	 	when 1000001101=> 
 	 	 	 	 <= C51515
 	 	 	when 1000001110=> 
 	 	 	 	 <= 760D0D
 	 	 	when 1000001111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1000010000=> 
 	 	 	 	 <= 7F0E0E
 	 	 	when 1000010001=> 
 	 	 	 	 <= C51515
 	 	 	when 1000010010=> 
 	 	 	 	 <= C51515
 	 	 	when 1000010011=> 
 	 	 	 	 <= C51515
 	 	 	when 1000010100=> 
 	 	 	 	 <= C51515
 	 	 	when 1000010101=> 
 	 	 	 	 <= C51515
 	 	 	when 1000010110=> 
 	 	 	 	 <= C51515
 	 	 	when 1000010111=> 
 	 	 	 	 <= C51515
 	 	 	when 1000011000=> 
 	 	 	 	 <= C51515
 	 	 	when 1000011001=> 
 	 	 	 	 <= C41414
 	 	 	when 1000011010=> 
 	 	 	 	 <= 810E0E
 	 	 	when 1000011011=> 
 	 	 	 	 <= 670B09
 	 	 	when 1000011100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1000011101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1000011110=> 
 	 	 	 	 <= 8C0G0G
 	 	 	when 1000100000=> 
 	 	 	 	 <= D74G4G
 	 	 	when 1000100001=> 
 	 	 	 	 <= C51515
 	 	 	when 1000100010=> 
 	 	 	 	 <= C41414
 	 	 	when 1000100011=> 
 	 	 	 	 <= BD1313
 	 	 	when 1000100100=> 
 	 	 	 	 <= 770D0D
 	 	 	when 1000100101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1000100110=> 
 	 	 	 	 <= B31212
 	 	 	when 1000100111=> 
 	 	 	 	 <= 9C1111
 	 	 	when 1000101000=> 
 	 	 	 	 <= 680B09
 	 	 	when 1000101001=> 
 	 	 	 	 <= 6B0B0B
 	 	 	when 1000101010=> 
 	 	 	 	 <= B81313
 	 	 	when 1000101011=> 
 	 	 	 	 <= C51515
 	 	 	when 1000101100=> 
 	 	 	 	 <= C51515
 	 	 	when 1000101101=> 
 	 	 	 	 <= C51515
 	 	 	when 1000101110=> 
 	 	 	 	 <= 7F0E0E
 	 	 	when 1000101111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1000110000=> 
 	 	 	 	 <= 750C0C
 	 	 	when 1000110001=> 
 	 	 	 	 <= C51515
 	 	 	when 1000110010=> 
 	 	 	 	 <= C51515
 	 	 	when 1000110011=> 
 	 	 	 	 <= C51515
 	 	 	when 1000110100=> 
 	 	 	 	 <= C51515
 	 	 	when 1000110101=> 
 	 	 	 	 <= C51515
 	 	 	when 1000110110=> 
 	 	 	 	 <= C51515
 	 	 	when 1000110111=> 
 	 	 	 	 <= C51515
 	 	 	when 1000111000=> 
 	 	 	 	 <= C11414
 	 	 	when 1000111001=> 
 	 	 	 	 <= 800E0E
 	 	 	when 1000111010=> 
 	 	 	 	 <= 67090B
 	 	 	when 1000111011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1000111100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1000111101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1000111110=> 
 	 	 	 	 <= 880F0F
 	 	 	when 1001000000=> 
 	 	 	 	 <= E47878
 	 	 	when 1001000001=> 
 	 	 	 	 <= C51515
 	 	 	when 1001000010=> 
 	 	 	 	 <= C51515
 	 	 	when 1001000011=> 
 	 	 	 	 <= C51515
 	 	 	when 1001000100=> 
 	 	 	 	 <= 910G0G
 	 	 	when 1001000101=> 
 	 	 	 	 <= 790D0D
 	 	 	when 1001000110=> 
 	 	 	 	 <= C01414
 	 	 	when 1001000111=> 
 	 	 	 	 <= C51515
 	 	 	when 1001001000=> 
 	 	 	 	 <= BC1313
 	 	 	when 1001001001=> 
 	 	 	 	 <= C01414
 	 	 	when 1001001010=> 
 	 	 	 	 <= C51515
 	 	 	when 1001001011=> 
 	 	 	 	 <= C51515
 	 	 	when 1001001100=> 
 	 	 	 	 <= C51515
 	 	 	when 1001001101=> 
 	 	 	 	 <= C31414
 	 	 	when 1001001110=> 
 	 	 	 	 <= 6E0B0B
 	 	 	when 1001001111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1001010000=> 
 	 	 	 	 <= 6D0B0B
 	 	 	when 1001010001=> 
 	 	 	 	 <= C41414
 	 	 	when 1001010010=> 
 	 	 	 	 <= C51515
 	 	 	when 1001010011=> 
 	 	 	 	 <= C51515
 	 	 	when 1001010100=> 
 	 	 	 	 <= C51515
 	 	 	when 1001010101=> 
 	 	 	 	 <= C51515
 	 	 	when 1001010110=> 
 	 	 	 	 <= C41414
 	 	 	when 1001010111=> 
 	 	 	 	 <= 9F1111
 	 	 	when 1001011000=> 
 	 	 	 	 <= 700C0C
 	 	 	when 1001011001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1001011010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1001011011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1001011100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1001011101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1001011110=> 
 	 	 	 	 <= 8C0G0G
 	 	 	when 1001100000=> 
 	 	 	 	 <= F7C5C5
 	 	 	when 1001100001=> 
 	 	 	 	 <= C51515
 	 	 	when 1001100010=> 
 	 	 	 	 <= C51515
 	 	 	when 1001100011=> 
 	 	 	 	 <= C51515
 	 	 	when 1001100100=> 
 	 	 	 	 <= C51515
 	 	 	when 1001100101=> 
 	 	 	 	 <= C51515
 	 	 	when 1001100110=> 
 	 	 	 	 <= C51515
 	 	 	when 1001100111=> 
 	 	 	 	 <= C51515
 	 	 	when 1001101000=> 
 	 	 	 	 <= C51515
 	 	 	when 1001101001=> 
 	 	 	 	 <= C51515
 	 	 	when 1001101010=> 
 	 	 	 	 <= C51515
 	 	 	when 1001101011=> 
 	 	 	 	 <= C51515
 	 	 	when 1001101100=> 
 	 	 	 	 <= C51515
 	 	 	when 1001101101=> 
 	 	 	 	 <= 8E0G0G
 	 	 	when 1001101110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1001101111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1001110000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1001110001=> 
 	 	 	 	 <= 760D0D
 	 	 	when 1001110010=> 
 	 	 	 	 <= 9C1111
 	 	 	when 1001110011=> 
 	 	 	 	 <= B71313
 	 	 	when 1001110100=> 
 	 	 	 	 <= B01212
 	 	 	when 1001110101=> 
 	 	 	 	 <= 8D0G0G
 	 	 	when 1001110110=> 
 	 	 	 	 <= 720C0C
 	 	 	when 1001110111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1001111000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1001111001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1001111010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1001111011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1001111100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1001111101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1001111110=> 
 	 	 	 	 <= B12626
 	 	 	when 1010000000=> 
 	 	 	 	 <= GDG7G7
 	 	 	when 1010000001=> 
 	 	 	 	 <= C61C1C
 	 	 	when 1010000010=> 
 	 	 	 	 <= C51515
 	 	 	when 1010000011=> 
 	 	 	 	 <= C51515
 	 	 	when 1010000100=> 
 	 	 	 	 <= C51515
 	 	 	when 1010000101=> 
 	 	 	 	 <= C51515
 	 	 	when 1010000110=> 
 	 	 	 	 <= C51515
 	 	 	when 1010000111=> 
 	 	 	 	 <= C51515
 	 	 	when 1010001000=> 
 	 	 	 	 <= C51515
 	 	 	when 1010001001=> 
 	 	 	 	 <= C51515
 	 	 	when 1010001010=> 
 	 	 	 	 <= C51515
 	 	 	when 1010001011=> 
 	 	 	 	 <= C41515
 	 	 	when 1010001100=> 
 	 	 	 	 <= 9E1111
 	 	 	when 1010001101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010001110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010001111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010010000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010010001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010010010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010010011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010010100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010010101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010010110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010010111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010011000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010011001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010011010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010011011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010011100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010011101=> 
 	 	 	 	 <= 6C0B0B
 	 	 	when 1010011110=> 
 	 	 	 	 <= E27979
 	 	 	when 1010100001=> 
 	 	 	 	 <= E17070
 	 	 	when 1010100010=> 
 	 	 	 	 <= C51515
 	 	 	when 1010100011=> 
 	 	 	 	 <= C51515
 	 	 	when 1010100100=> 
 	 	 	 	 <= C51515
 	 	 	when 1010100101=> 
 	 	 	 	 <= C51515
 	 	 	when 1010100110=> 
 	 	 	 	 <= C51515
 	 	 	when 1010100111=> 
 	 	 	 	 <= C51515
 	 	 	when 1010101000=> 
 	 	 	 	 <= C51515
 	 	 	when 1010101001=> 
 	 	 	 	 <= C51415
 	 	 	when 1010101010=> 
 	 	 	 	 <= C11414
 	 	 	when 1010101011=> 
 	 	 	 	 <= 8D0G0G
 	 	 	when 1010101100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010101101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010101110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010101111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010110000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010110001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010110010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010110011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010110100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010110101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010110110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010110111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010111000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010111001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010111010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010111011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010111100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1010111101=> 
 	 	 	 	 <= 921010
 	 	 	when 1010111110=> 
 	 	 	 	 <= G4EEEE
 	 	 	when 1011000001=> 
 	 	 	 	 <= G6F4F4
 	 	 	when 1011000010=> 
 	 	 	 	 <= C61818
 	 	 	when 1011000011=> 
 	 	 	 	 <= C51515
 	 	 	when 1011000100=> 
 	 	 	 	 <= C51515
 	 	 	when 1011000101=> 
 	 	 	 	 <= C51515
 	 	 	when 1011000110=> 
 	 	 	 	 <= C51515
 	 	 	when 1011000111=> 
 	 	 	 	 <= C41415
 	 	 	when 1011001000=> 
 	 	 	 	 <= B31212
 	 	 	when 1011001001=> 
 	 	 	 	 <= 7F0E0E
 	 	 	when 1011001010=> 
 	 	 	 	 <= 690B0B
 	 	 	when 1011001011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011001100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011001101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011001110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011001111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011010000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011010001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011010010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011010011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011010100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011010101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011010110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011010111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011011000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011011001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011011010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011011011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011011100=> 
 	 	 	 	 <= 710C0C
 	 	 	when 1011011101=> 
 	 	 	 	 <= DD6363
 	 	 	when 1011100010=> 
 	 	 	 	 <= E98889
 	 	 	when 1011100011=> 
 	 	 	 	 <= C51515
 	 	 	when 1011100100=> 
 	 	 	 	 <= C51515
 	 	 	when 1011100101=> 
 	 	 	 	 <= C51515
 	 	 	when 1011100110=> 
 	 	 	 	 <= C41414
 	 	 	when 1011100111=> 
 	 	 	 	 <= 810E0E
 	 	 	when 1011101000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011101001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011101010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011101011=> 
 	 	 	 	 <= 7E0E0E
 	 	 	when 1011101100=> 
 	 	 	 	 <= 941010
 	 	 	when 1011101101=> 
 	 	 	 	 <= 910G10
 	 	 	when 1011101110=> 
 	 	 	 	 <= 730C0C
 	 	 	when 1011101111=> 
 	 	 	 	 <= 680B09
 	 	 	when 1011110000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011110001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011110010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011110011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011110100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011110101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011110110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011110111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011111000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011111001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011111010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1011111011=> 
 	 	 	 	 <= 6C0B0B
 	 	 	when 1011111100=> 
 	 	 	 	 <= BB1E1E
 	 	 	when 1011111101=> 
 	 	 	 	 <= G8F9F9
 	 	 	when 1100000010=> 
 	 	 	 	 <= GFGDGD
 	 	 	when 1100000011=> 
 	 	 	 	 <= D54848
 	 	 	when 1100000100=> 
 	 	 	 	 <= C51515
 	 	 	when 1100000101=> 
 	 	 	 	 <= C51515
 	 	 	when 1100000110=> 
 	 	 	 	 <= 8G0G0G
 	 	 	when 1100000111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100001000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100001001=> 
 	 	 	 	 <= 8B0F0F
 	 	 	when 1100001010=> 
 	 	 	 	 <= BD1313
 	 	 	when 1100001011=> 
 	 	 	 	 <= C51414
 	 	 	when 1100001100=> 
 	 	 	 	 <= C51515
 	 	 	when 1100001101=> 
 	 	 	 	 <= C51515
 	 	 	when 1100001110=> 
 	 	 	 	 <= C41414
 	 	 	when 1100001111=> 
 	 	 	 	 <= 9F1111
 	 	 	when 1100010000=> 
 	 	 	 	 <= 6D0B0B
 	 	 	when 1100010001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100010010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100010011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100010100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100010101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100010110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100010111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100011000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100011001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100011010=> 
 	 	 	 	 <= 690B0B
 	 	 	when 1100011011=> 
 	 	 	 	 <= B31212
 	 	 	when 1100011100=> 
 	 	 	 	 <= F6C0C0
 	 	 	when 1100100011=> 
 	 	 	 	 <= G9FGFG
 	 	 	when 1100100100=> 
 	 	 	 	 <= CG3535
 	 	 	when 1100100101=> 
 	 	 	 	 <= C51515
 	 	 	when 1100100110=> 
 	 	 	 	 <= 740C0C
 	 	 	when 1100100111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100101000=> 
 	 	 	 	 <= 910G0G
 	 	 	when 1100101001=> 
 	 	 	 	 <= C41515
 	 	 	when 1100101010=> 
 	 	 	 	 <= C51515
 	 	 	when 1100101011=> 
 	 	 	 	 <= C51515
 	 	 	when 1100101100=> 
 	 	 	 	 <= C51515
 	 	 	when 1100101101=> 
 	 	 	 	 <= C51515
 	 	 	when 1100101110=> 
 	 	 	 	 <= C51515
 	 	 	when 1100101111=> 
 	 	 	 	 <= C51515
 	 	 	when 1100110000=> 
 	 	 	 	 <= B41212
 	 	 	when 1100110001=> 
 	 	 	 	 <= 690B0B
 	 	 	when 1100110010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100110011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100110100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100110101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100110110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100110111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100111000=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1100111001=> 
 	 	 	 	 <= 6B0B0B
 	 	 	when 1100111010=> 
 	 	 	 	 <= B01112
 	 	 	when 1100111011=> 
 	 	 	 	 <= EC8F8F
 	 	 	when 1101000100=> 
 	 	 	 	 <= G9FEFE
 	 	 	when 1101000101=> 
 	 	 	 	 <= D24040
 	 	 	when 1101000110=> 
 	 	 	 	 <= B01212
 	 	 	when 1101000111=> 
 	 	 	 	 <= 92100G
 	 	 	when 1101001000=> 
 	 	 	 	 <= C41414
 	 	 	when 1101001001=> 
 	 	 	 	 <= C51515
 	 	 	when 1101001010=> 
 	 	 	 	 <= C51515
 	 	 	when 1101001011=> 
 	 	 	 	 <= C51515
 	 	 	when 1101001100=> 
 	 	 	 	 <= C51515
 	 	 	when 1101001101=> 
 	 	 	 	 <= C51515
 	 	 	when 1101001110=> 
 	 	 	 	 <= C51515
 	 	 	when 1101001111=> 
 	 	 	 	 <= C51515
 	 	 	when 1101010000=> 
 	 	 	 	 <= C51515
 	 	 	when 1101010001=> 
 	 	 	 	 <= 921010
 	 	 	when 1101010010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1101010011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1101010100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1101010101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1101010110=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1101010111=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1101011000=> 
 	 	 	 	 <= 6G0C0C
 	 	 	when 1101011001=> 
 	 	 	 	 <= B61313
 	 	 	when 1101011010=> 
 	 	 	 	 <= EE9494
 	 	 	when 1101100101=> 
 	 	 	 	 <= GEG9G9
 	 	 	when 1101100110=> 
 	 	 	 	 <= E27373
 	 	 	when 1101100111=> 
 	 	 	 	 <= C51515
 	 	 	when 1101101000=> 
 	 	 	 	 <= C51515
 	 	 	when 1101101001=> 
 	 	 	 	 <= C51515
 	 	 	when 1101101010=> 
 	 	 	 	 <= C51515
 	 	 	when 1101101011=> 
 	 	 	 	 <= C51515
 	 	 	when 1101101100=> 
 	 	 	 	 <= C51515
 	 	 	when 1101101101=> 
 	 	 	 	 <= C51515
 	 	 	when 1101101110=> 
 	 	 	 	 <= C51515
 	 	 	when 1101101111=> 
 	 	 	 	 <= C51515
 	 	 	when 1101110000=> 
 	 	 	 	 <= C41515
 	 	 	when 1101110001=> 
 	 	 	 	 <= 951010
 	 	 	when 1101110010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1101110011=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1101110100=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1101110101=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1101110110=> 
 	 	 	 	 <= 690B0B
 	 	 	when 1101110111=> 
 	 	 	 	 <= 8C0G0G
 	 	 	when 1101111000=> 
 	 	 	 	 <= C82828
 	 	 	when 1101111001=> 
 	 	 	 	 <= FCD0D0
 	 	 	when 1110000110=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1110000111=> 
 	 	 	 	 <= FGDEDE
 	 	 	when 1110001000=> 
 	 	 	 	 <= D44747
 	 	 	when 1110001001=> 
 	 	 	 	 <= C41415
 	 	 	when 1110001010=> 
 	 	 	 	 <= C51515
 	 	 	when 1110001011=> 
 	 	 	 	 <= C51515
 	 	 	when 1110001100=> 
 	 	 	 	 <= C51515
 	 	 	when 1110001101=> 
 	 	 	 	 <= C51515
 	 	 	when 1110001110=> 
 	 	 	 	 <= C51515
 	 	 	when 1110001111=> 
 	 	 	 	 <= C51515
 	 	 	when 1110010000=> 
 	 	 	 	 <= BB1313
 	 	 	when 1110010001=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1110010010=> 
 	 	 	 	 <= 680B0B
 	 	 	when 1110010011=> 
 	 	 	 	 <= 680B09
 	 	 	when 1110010100=> 
 	 	 	 	 <= 6D0B0B
 	 	 	when 1110010101=> 
 	 	 	 	 <= 8B0F0F
 	 	 	when 1110010110=> 
 	 	 	 	 <= C11B1B
 	 	 	when 1110010111=> 
 	 	 	 	 <= E67G7G
 	 	 	when 1110011000=> 
 	 	 	 	 <= GCG4G4
 	 	 	when 1110101000=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1110101001=> 
 	 	 	 	 <= FGDGDG
 	 	 	when 1110101010=> 
 	 	 	 	 <= E27070
 	 	 	when 1110101011=> 
 	 	 	 	 <= CB2727
 	 	 	when 1110101100=> 
 	 	 	 	 <= C41415
 	 	 	when 1110101101=> 
 	 	 	 	 <= C41515
 	 	 	when 1110101110=> 
 	 	 	 	 <= C51515
 	 	 	when 1110101111=> 
 	 	 	 	 <= C51515
 	 	 	when 1110110000=> 
 	 	 	 	 <= C31414
 	 	 	when 1110110001=> 
 	 	 	 	 <= 880F0F
 	 	 	when 1110110010=> 
 	 	 	 	 <= 880F0F
 	 	 	when 1110110011=> 
 	 	 	 	 <= 9E1212
 	 	 	when 1110110100=> 
 	 	 	 	 <= D24445
 	 	 	when 1110110101=> 
 	 	 	 	 <= EF9898
 	 	 	when 1110110110=> 
 	 	 	 	 <= GBG1G1
 	 	 	when 1111001011=> 
 	 	 	 	 <= GFGFGF
 	 	 	when 1111001100=> 
 	 	 	 	 <= G6F3F3
 	 	 	when 1111001101=> 
 	 	 	 	 <= F9CBCB
 	 	 	when 1111001110=> 
 	 	 	 	 <= F09F9F
 	 	 	when 1111001111=> 
 	 	 	 	 <= EE9494
 	 	 	when 1111010000=> 
 	 	 	 	 <= EF9797
 	 	 	when 1111010001=> 
 	 	 	 	 <= F3B8B8
 	 	 	when 1111010010=> 
 	 	 	 	 <= FFDBDB
 	 	 	when 1111010011=> 
 	 	 	 	 <= GDG6G6
 	 	 	when 1111010100=> 
 	 	 	 	 <= GFGFGF 
 	 	 end case; 
     	 end if;  
     end process; 
 address <= row & col; 
 end;
